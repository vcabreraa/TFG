------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : mri1_256x256.pgm 
--- Filas    : 256 
--- Columnas : 256 
--- Color    :  8 bits



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 8 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;

library WORK;
use WORK.IMG_PKG.ALL; 

library WORK;
use WORK.IMG_PKG.ALL; 


entity R1sp is
  port (
    clk  : in  std_logic;   -- reloj    
    addr1 : in  std_logic_vector(c_2dim_img-1 downto 0);
    dout1 : out std_logic_vector(8-1 downto 0) 
  );
end R1sp;


architecture BEHAVIORAL of R1sp is
  
  signal addr1_int  : natural range 0 to 2**c_2dim_img-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant filaimg : memostruct := (
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010100",
       "00001010",
       "00010111",
       "00100000",
       "00011110",
       "00010011",
       "00001101",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001000",
       "00000111",
       "00001100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001111",
       "00011110",
       "00110001",
       "00110100",
       "00110010",
       "00101001",
       "00010001",
       "00001101",
       "00010010",
       "00001000",
       "00001010",
       "00001111",
       "00011010",
       "00100011",
       "00011011",
       "00001111",
       "00001010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00110010",
       "00111011",
       "00101111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001101",
       "00011000",
       "00010111",
       "00010110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001101",
       "00011101",
       "00111000",
       "00110100",
       "00110100",
       "00110001",
       "00110101",
       "00100101",
       "00001100",
       "00001111",
       "00001000",
       "00010001",
       "00101010",
       "00110010",
       "00110001",
       "00101001",
       "00011101",
       "00010001",
       "00001001",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00110001",
       "00111000",
       "00000000",
       "00000000",
       "00000000",
       "00111111",
       "00111110",
       "00110011",
       "00110010",
       "00110001",
       "00010101",
       "00011000",
       "00011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010001",
       "00100001",
       "00101111",
       "00101010",
       "00101000",
       "00011101",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001011",
       "00110011",
       "00110101",
       "00101111",
       "00110010",
       "00101111",
       "00110010",
       "00110001",
       "00011000",
       "00001001",
       "00001010",
       "00100101",
       "00110011",
       "00110001",
       "00110000",
       "00110001",
       "00101101",
       "00011100",
       "00010001",
       "00001110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00110110",
       "00111011",
       "00110100",
       "00000000",
       "00000000",
       "00110110",
       "00101111",
       "00101110",
       "00100110",
       "00011101",
       "00011101",
       "00010100",
       "00010110",
       "00010101",
       "00001010",
       "00001011",
       "00001100",
       "00001011",
       "00001001",
       "00001000",
       "00100001",
       "00101111",
       "00110001",
       "00101110",
       "00110010",
       "00101100",
       "00001111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010100",
       "00111000",
       "00101111",
       "00111000",
       "00110111",
       "00111001",
       "00110001",
       "00110011",
       "00100111",
       "00001101",
       "00010010",
       "00110100",
       "00101101",
       "00101111",
       "00101110",
       "00110011",
       "00110101",
       "00100110",
       "00010000",
       "00010011",
       "00010011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00111011",
       "00110001",
       "00110110",
       "00110100",
       "00111000",
       "00111001",
       "00101100",
       "00011100",
       "00010101",
       "00101110",
       "00101111",
       "00101101",
       "00100101",
       "00011111",
       "00010110",
       "00001111",
       "00001001",
       "00001010",
       "00001011",
       "00000110",
       "00010011",
       "00110000",
       "00101110",
       "00110000",
       "00101101",
       "00110001",
       "00110000",
       "00011110",
       "00000101",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00011100",
       "00011010",
       "00110010",
       "00101110",
       "00111100",
       "00111111",
       "01000001",
       "00110111",
       "00110100",
       "00101111",
       "00010110",
       "00011101",
       "00110110",
       "00110001",
       "00111011",
       "00111001",
       "00110000",
       "00110001",
       "00100110",
       "00011111",
       "00101000",
       "00100011",
       "00011101",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00111100",
       "00111001",
       "00101111",
       "00110101",
       "00101111",
       "00111101",
       "00110001",
       "00010101",
       "00010110",
       "00101101",
       "00111001",
       "00110000",
       "00101111",
       "00101111",
       "00110000",
       "00101100",
       "00011100",
       "00000111",
       "00001010",
       "00001000",
       "00001010",
       "00100100",
       "00110111",
       "00101111",
       "00110101",
       "00101111",
       "00101111",
       "00101101",
       "00101011",
       "00001001",
       "00001011",
       "00000011",
       "00010001",
       "00001000",
       "00011100",
       "00011111",
       "00011000",
       "00110011",
       "00101101",
       "00111011",
       "01000010",
       "01000110",
       "00111110",
       "00110100",
       "00101111",
       "00100001",
       "00100000",
       "00110100",
       "00110101",
       "01000011",
       "00111111",
       "00110011",
       "00110000",
       "00100011",
       "00101011",
       "00110100",
       "00110000",
       "00101111",
       "00100111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "01000111",
       "00111001",
       "00111001",
       "00110001",
       "00111011",
       "00111111",
       "00011110",
       "00010010",
       "00001101",
       "00011111",
       "00110110",
       "00101111",
       "00101101",
       "00110011",
       "00101100",
       "00110000",
       "00110101",
       "00110001",
       "00001111",
       "00000111",
       "00000101",
       "00010010",
       "00101111",
       "00110110",
       "00110110",
       "00111010",
       "00110111",
       "00110011",
       "00101110",
       "00110001",
       "00010111",
       "00001001",
       "00000111",
       "00010100",
       "00000111",
       "00011101",
       "00100001",
       "00010001",
       "00110011",
       "00101111",
       "00110110",
       "00111111",
       "01001000",
       "01000001",
       "00111001",
       "00101111",
       "00101001",
       "00100010",
       "00110001",
       "00110110",
       "01000100",
       "00111100",
       "00110101",
       "00101010",
       "00100111",
       "00110001",
       "00110100",
       "00110111",
       "00110100",
       "00110010",
       "00100111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00111011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00111010",
       "00110001",
       "00100100",
       "00101111",
       "00111011",
       "00110011",
       "00011000",
       "00001010",
       "00010001",
       "00001101",
       "00100000",
       "00110011",
       "00110010",
       "00110100",
       "00111101",
       "00110110",
       "00110010",
       "00101100",
       "00110110",
       "00100001",
       "00000111",
       "00000101",
       "00011110",
       "00110010",
       "00110001",
       "00111000",
       "01000000",
       "01000010",
       "00111000",
       "00110000",
       "00110010",
       "00100111",
       "00001001",
       "00001100",
       "00011011",
       "00000110",
       "00011111",
       "00100010",
       "00001100",
       "00101001",
       "00101110",
       "00110010",
       "00110101",
       "01000010",
       "01000001",
       "00111100",
       "00110011",
       "00101100",
       "00101001",
       "00110000",
       "00111011",
       "01000110",
       "00111001",
       "00110001",
       "00100100",
       "00101101",
       "00110101",
       "00110010",
       "00110100",
       "00110101",
       "00110101",
       "00110001",
       "00011010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00110110",
       "00110100",
       "00111110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00011100",
       "00011010",
       "00100010",
       "00110010",
       "00011111",
       "00011000",
       "00011001",
       "00010100",
       "00001001",
       "00000111",
       "00100000",
       "00110111",
       "00101111",
       "00110100",
       "01000100",
       "01000010",
       "00111010",
       "00110011",
       "00110101",
       "00110010",
       "00001111",
       "00000110",
       "00100110",
       "00110001",
       "00110011",
       "00111010",
       "01000101",
       "01000101",
       "00111100",
       "00110000",
       "00110001",
       "00101001",
       "00010000",
       "00010101",
       "00011001",
       "00000111",
       "00100001",
       "00100111",
       "00000111",
       "00011110",
       "00101011",
       "00110101",
       "00101101",
       "00111100",
       "01000001",
       "01000011",
       "00111110",
       "00110001",
       "00101110",
       "00110010",
       "01000000",
       "01000100",
       "00110101",
       "00101100",
       "00101011",
       "00111010",
       "00110110",
       "00110011",
       "00110101",
       "00110110",
       "00110010",
       "00110011",
       "00011100",
       "00000000",
       "00000000",
       "00000111",
       "00001100",
       "00010110",
       "00001111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00110100",
       "00110010",
       "00110110",
       "00101110",
       "00110101",
       "00110100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010111",
       "00010011",
       "00010000",
       "00100011",
       "00011101",
       "00100100",
       "00101001",
       "00101101",
       "00101000",
       "00011000",
       "00001011",
       "00001000",
       "00010110",
       "00101110",
       "00110001",
       "00110100",
       "00111111",
       "01000111",
       "01000011",
       "00111101",
       "00110000",
       "00110101",
       "00010111",
       "00000111",
       "00101110",
       "00101101",
       "00110101",
       "00111101",
       "01000101",
       "00111111",
       "00111010",
       "00110010",
       "00110100",
       "00101000",
       "00011001",
       "00011111",
       "00010010",
       "00001000",
       "00100101",
       "00101001",
       "00000100",
       "00001101",
       "00100000",
       "00110101",
       "00101111",
       "00110101",
       "00111011",
       "01001010",
       "01000111",
       "00111110",
       "00110101",
       "00111011",
       "01000101",
       "01000011",
       "00110011",
       "00101100",
       "00110011",
       "00110101",
       "00110101",
       "00110110",
       "00110101",
       "00110100",
       "00110011",
       "00110001",
       "00011010",
       "00001001",
       "00001001",
       "00001110",
       "00001111",
       "00011101",
       "00101000",
       "00010010",
       "00100000",
       "00000000",
       "00101111",
       "00110100",
       "00110110",
       "00101110",
       "00101100",
       "00110000",
       "00110011",
       "00101100",
       "00010111",
       "01110011",
       "10111100",
       "10100101",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010100",
       "00011001",
       "00100010",
       "00010110",
       "00011010",
       "00101111",
       "00111101",
       "00110110",
       "00110001",
       "00100110",
       "00010110",
       "00001010",
       "00010011",
       "00101101",
       "00110110",
       "00110100",
       "00111011",
       "01000011",
       "01000101",
       "01000100",
       "00110011",
       "00110011",
       "00100010",
       "00001101",
       "00110010",
       "00101100",
       "00111101",
       "01000011",
       "01000101",
       "00111011",
       "00110111",
       "00110011",
       "00110010",
       "00100100",
       "00100100",
       "00011101",
       "00010000",
       "00000111",
       "00100010",
       "00101000",
       "00000100",
       "00000110",
       "00001011",
       "00100011",
       "00101011",
       "00110101",
       "00101111",
       "01000000",
       "01000110",
       "01000110",
       "01000110",
       "01001001",
       "01000110",
       "01000011",
       "00101111",
       "00101111",
       "00110101",
       "00110010",
       "00110111",
       "00110111",
       "00110110",
       "00110101",
       "00110101",
       "00100111",
       "00010010",
       "00001001",
       "00001010",
       "00001010",
       "00010011",
       "00101111",
       "00110110",
       "01000010",
       "00101100",
       "00010101",
       "00110101",
       "00111011",
       "01001001",
       "00111111",
       "01000010",
       "00110100",
       "00101101",
       "00111011",
       "00110000",
       "00100001",
       "01010010",
       "10111001",
       "10110111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010010",
       "00011111",
       "00101001",
       "00011011",
       "00011111",
       "00110101",
       "00110101",
       "00110001",
       "00110110",
       "00110101",
       "00101001",
       "00011001",
       "00001011",
       "00010001",
       "00101110",
       "00110101",
       "00110011",
       "00111000",
       "01000011",
       "01001001",
       "01000111",
       "00111010",
       "00110001",
       "00101001",
       "00011100",
       "00110011",
       "00110010",
       "01001010",
       "01000100",
       "01000111",
       "00110100",
       "00101111",
       "00101100",
       "00101001",
       "00100010",
       "00101100",
       "00011110",
       "00010011",
       "00000111",
       "00100001",
       "00101001",
       "00000101",
       "00001110",
       "00001001",
       "00010100",
       "00010111",
       "00101111",
       "00101111",
       "00110101",
       "01000011",
       "01001001",
       "01001101",
       "01001110",
       "01000111",
       "01000011",
       "00110010",
       "00110100",
       "00111010",
       "00111101",
       "00111100",
       "00111001",
       "00111000",
       "00110111",
       "00110010",
       "00011111",
       "00001100",
       "00001010",
       "00001001",
       "00001111",
       "00100110",
       "00111001",
       "00110101",
       "00110100",
       "00111100",
       "00101111",
       "00010100",
       "00111100",
       "00110101",
       "00111101",
       "01001110",
       "01000100",
       "00111010",
       "00111001",
       "00111110",
       "00101100",
       "00111011",
       "01000001",
       "11000011",
       "10100111",
       "10011001",
       "10000110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00011111",
       "00011011",
       "00010101",
       "00100111",
       "00111010",
       "00110001",
       "00110001",
       "00110111",
       "00110111",
       "00110100",
       "00110000",
       "00011111",
       "00010000",
       "00010000",
       "00101001",
       "00110011",
       "00110001",
       "00111001",
       "01000110",
       "01001001",
       "01001001",
       "01000001",
       "00110101",
       "00101100",
       "00101101",
       "00110101",
       "00111010",
       "01001101",
       "01000110",
       "01000000",
       "00101111",
       "00101101",
       "00101000",
       "00101100",
       "00101110",
       "00110011",
       "00100011",
       "00011011",
       "00000101",
       "00100010",
       "00101010",
       "00000100",
       "00010001",
       "00001100",
       "00010100",
       "00001100",
       "00010100",
       "00100110",
       "00110100",
       "00111100",
       "01001000",
       "01001001",
       "01001101",
       "01001101",
       "01000111",
       "00111111",
       "00111111",
       "01000100",
       "01000111",
       "01000000",
       "00111011",
       "00110100",
       "00110110",
       "00101101",
       "00011011",
       "00001101",
       "00001101",
       "00000110",
       "00010100",
       "00110110",
       "00111010",
       "00110111",
       "00111001",
       "00110000",
       "00111010",
       "00101000",
       "00001001",
       "00101010",
       "00101101",
       "00111010",
       "01000010",
       "00111001",
       "00111011",
       "01000101",
       "01000101",
       "00101100",
       "00101111",
       "01000110",
       "10111100",
       "10101001",
       "01111110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00110011",
       "00100100",
       "00010111",
       "00101010",
       "00110110",
       "00101110",
       "00110000",
       "00111100",
       "00111101",
       "00111001",
       "00111001",
       "00110100",
       "00100010",
       "00010011",
       "00010011",
       "00101011",
       "00110100",
       "00110110",
       "00111101",
       "01000110",
       "01001001",
       "01001100",
       "01001000",
       "00111100",
       "00110000",
       "00110001",
       "00110111",
       "01000101",
       "01001100",
       "01001000",
       "00111001",
       "00101111",
       "00101100",
       "00101101",
       "00110011",
       "00110001",
       "00111000",
       "00101111",
       "00101100",
       "00001010",
       "00011011",
       "00101010",
       "00000011",
       "00001101",
       "00001011",
       "00010101",
       "00010001",
       "00001010",
       "00010001",
       "00101010",
       "00110101",
       "01000010",
       "01001110",
       "01001111",
       "01001101",
       "01001101",
       "01001011",
       "01001100",
       "01001101",
       "01001100",
       "01000000",
       "00111001",
       "00110011",
       "00110111",
       "00101001",
       "00010110",
       "00001110",
       "00001100",
       "00000111",
       "00100101",
       "00111010",
       "00111010",
       "01000110",
       "01000100",
       "00111011",
       "00110010",
       "00101101",
       "00010101",
       "00000101",
       "00100110",
       "00100010",
       "01000101",
       "01000110",
       "01000000",
       "01000000",
       "00111011",
       "00111111",
       "00101001",
       "00100010",
       "01001001",
       "10101100",
       "10010100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00100100",
       "00011000",
       "00110101",
       "00110110",
       "00110000",
       "00110100",
       "00111010",
       "01000010",
       "01001010",
       "00111111",
       "00110110",
       "00110000",
       "00100111",
       "00011001",
       "00010100",
       "00101101",
       "00111001",
       "00111001",
       "00111101",
       "01000110",
       "01010001",
       "01001100",
       "01001111",
       "01000100",
       "00111010",
       "00111000",
       "01000010",
       "01001100",
       "01001010",
       "01000100",
       "00111000",
       "00101111",
       "00101110",
       "00101111",
       "00110101",
       "00110001",
       "00111000",
       "00110010",
       "00110101",
       "00010001",
       "00010110",
       "00100100",
       "00000100",
       "00001011",
       "00001011",
       "00001111",
       "00001110",
       "00010010",
       "00011001",
       "00101000",
       "00110011",
       "00111110",
       "01001110",
       "01001110",
       "01001101",
       "01001111",
       "01010100",
       "01010001",
       "01001110",
       "01001011",
       "01000001",
       "00110111",
       "00110100",
       "00110110",
       "00100001",
       "00001111",
       "00001011",
       "00001011",
       "00010001",
       "00110101",
       "00111110",
       "01000100",
       "01001011",
       "00111111",
       "00111000",
       "00110111",
       "00100011",
       "00001100",
       "00001010",
       "00010001",
       "00100110",
       "00111101",
       "00111001",
       "00111101",
       "00111110",
       "00101111",
       "00110100",
       "00110101",
       "00100101",
       "00101101",
       "00111000",
       "10110010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00011110",
       "00011000",
       "00101111",
       "00110101",
       "00101100",
       "00110110",
       "00110110",
       "01000011",
       "01000110",
       "01000111",
       "00111101",
       "00111010",
       "00110100",
       "00110010",
       "00011010",
       "00010100",
       "00101100",
       "00111000",
       "00111000",
       "01000001",
       "01000111",
       "01001111",
       "01001110",
       "01010010",
       "01001100",
       "01001100",
       "01001011",
       "01001100",
       "01001101",
       "01001001",
       "00111101",
       "00110011",
       "00101111",
       "00110001",
       "00110001",
       "00110010",
       "00110101",
       "00110111",
       "00110010",
       "00110000",
       "00011001",
       "00010011",
       "00011001",
       "00000100",
       "00001100",
       "00001001",
       "00001100",
       "00001110",
       "00011011",
       "00101010",
       "00110100",
       "00110101",
       "00111110",
       "01001101",
       "01001110",
       "01001111",
       "01001111",
       "01010100",
       "01001111",
       "01001110",
       "01001010",
       "00111111",
       "00110111",
       "00110100",
       "00110010",
       "00011011",
       "00001010",
       "00001010",
       "00001100",
       "00101101",
       "00110111",
       "00111111",
       "01001110",
       "01000011",
       "00111000",
       "00110011",
       "00100111",
       "00011111",
       "00001011",
       "00001010",
       "00001111",
       "00011110",
       "00101000",
       "00110111",
       "00110001",
       "00111100",
       "01000001",
       "00111000",
       "00110111",
       "00101100",
       "00100111",
       "00101011",
       "01010110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010100",
       "00010101",
       "00110100",
       "00110001",
       "00110010",
       "00110111",
       "00110111",
       "00111101",
       "01000111",
       "01000111",
       "01001001",
       "01000101",
       "00111001",
       "00110111",
       "00110011",
       "00100011",
       "00011001",
       "00101110",
       "00111001",
       "00111011",
       "01000000",
       "01001101",
       "01001111",
       "01001111",
       "01001100",
       "01001111",
       "01001111",
       "01001100",
       "01001001",
       "01001001",
       "01001000",
       "00110111",
       "00101110",
       "00110001",
       "00110000",
       "00110011",
       "00110010",
       "00110101",
       "00111000",
       "00110011",
       "00110011",
       "00011011",
       "00001111",
       "00010110",
       "00001001",
       "00001100",
       "00001001",
       "00001101",
       "00001111",
       "00011100",
       "00101111",
       "00111010",
       "00111001",
       "01000001",
       "01001111",
       "01010101",
       "01010010",
       "01010010",
       "01010011",
       "01010010",
       "01010101",
       "01001011",
       "00111100",
       "00110011",
       "00110110",
       "00101111",
       "00010111",
       "00001010",
       "00001100",
       "00011111",
       "00111101",
       "00111001",
       "01001001",
       "01001001",
       "00111110",
       "00110100",
       "00100001",
       "00010111",
       "00010001",
       "00001100",
       "00001100",
       "00001110",
       "00011110",
       "00011011",
       "00101001",
       "00110001",
       "00111001",
       "01000100",
       "01000001",
       "00101110",
       "00101100",
       "00110010",
       "00101000",
       "00011010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010010",
       "00101111",
       "00110010",
       "00110100",
       "00110110",
       "00110101",
       "01000000",
       "00111110",
       "01000111",
       "01000111",
       "01001100",
       "01001001",
       "00111100",
       "00110110",
       "00110010",
       "00101110",
       "00011110",
       "00101100",
       "00111001",
       "00111010",
       "00111100",
       "01001000",
       "01010010",
       "01001111",
       "01010001",
       "01010011",
       "01001111",
       "01001101",
       "01001100",
       "01000111",
       "01000000",
       "00110101",
       "00101101",
       "00110011",
       "00110000",
       "00110111",
       "00110110",
       "00110100",
       "00110110",
       "00101101",
       "00110011",
       "00010111",
       "00001111",
       "00011101",
       "00001000",
       "00010010",
       "00001100",
       "00001111",
       "00001111",
       "00010110",
       "00101000",
       "00111011",
       "00110110",
       "01000010",
       "01001101",
       "01010001",
       "01010100",
       "01001111",
       "01010100",
       "01010001",
       "01010100",
       "01001100",
       "00111110",
       "00110110",
       "00111000",
       "00101000",
       "00010100",
       "00001011",
       "00011011",
       "00110101",
       "00111011",
       "01000000",
       "01001111",
       "01000000",
       "00111010",
       "00100101",
       "00001110",
       "00001011",
       "00001011",
       "00001010",
       "00001011",
       "00010011",
       "00001101",
       "00010101",
       "00001111",
       "00101010",
       "01001111",
       "00110011",
       "01001101",
       "00111010",
       "00101000",
       "00110100",
       "00111110",
       "00011101",
       "00101010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010100",
       "00101011",
       "00101110",
       "00110000",
       "00101110",
       "00110011",
       "00110110",
       "00111101",
       "00111101",
       "01000110",
       "01001001",
       "01001100",
       "01001100",
       "01000111",
       "00110110",
       "00110010",
       "00101100",
       "00011101",
       "00100101",
       "00111010",
       "00111010",
       "01000000",
       "01000001",
       "01001110",
       "01010000",
       "01010100",
       "01010101",
       "01010101",
       "01010010",
       "01001110",
       "01000110",
       "00111101",
       "00110010",
       "00110010",
       "00110010",
       "00101100",
       "00110110",
       "00110100",
       "00101110",
       "00110010",
       "00101011",
       "00101100",
       "00010011",
       "00010000",
       "00011111",
       "00001110",
       "00011000",
       "00010001",
       "00010000",
       "00010010",
       "00010100",
       "00100001",
       "00110100",
       "00110101",
       "01000001",
       "01001100",
       "01001011",
       "01010000",
       "01010000",
       "01010011",
       "01010011",
       "01010000",
       "01001001",
       "01000001",
       "00111010",
       "00111000",
       "00100000",
       "00001111",
       "00010001",
       "00110011",
       "00111010",
       "00111011",
       "01001001",
       "01010000",
       "00111110",
       "00110111",
       "00010110",
       "00001010",
       "00001001",
       "00001101",
       "00001111",
       "00001100",
       "00001110",
       "00010010",
       "00001100",
       "00010010",
       "00010110",
       "00110001",
       "00110101",
       "01000100",
       "01000100",
       "00101000",
       "00111110",
       "00110000",
       "00110011",
       "00100011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00110110",
       "00001110",
       "00101100",
       "00101101",
       "00110110",
       "00101111",
       "00101110",
       "00110001",
       "00110000",
       "00110011",
       "00111010",
       "01000010",
       "01000111",
       "01001110",
       "01010001",
       "01001100",
       "00111110",
       "00110111",
       "00101100",
       "00011000",
       "00011110",
       "00110110",
       "00110111",
       "01000111",
       "01000110",
       "01001000",
       "01010001",
       "01010011",
       "01010101",
       "01010100",
       "01010011",
       "01010001",
       "01000111",
       "00111001",
       "00110010",
       "00110011",
       "00110000",
       "00100101",
       "00101011",
       "00101011",
       "00100101",
       "00101011",
       "00100100",
       "00100001",
       "00001010",
       "00011000",
       "00100101",
       "00010010",
       "00011010",
       "00010011",
       "00010010",
       "00010011",
       "00001111",
       "00010111",
       "00100110",
       "00110110",
       "00111110",
       "01010000",
       "01001101",
       "01010011",
       "01010011",
       "01010110",
       "01011000",
       "01001111",
       "01001000",
       "00111111",
       "00111010",
       "00111000",
       "00011001",
       "00001010",
       "00101101",
       "00111001",
       "00111100",
       "01000111",
       "01010001",
       "01001010",
       "00111011",
       "00110101",
       "00010011",
       "00001101",
       "00001110",
       "00001100",
       "00000111",
       "00010000",
       "00001110",
       "00010010",
       "00001111",
       "00001110",
       "00010100",
       "00010011",
       "00011111",
       "00111011",
       "01000010",
       "00111000",
       "00110110",
       "00110000",
       "00110011",
       "00101001",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010111",
       "00011110",
       "00101111",
       "00110110",
       "00110000",
       "00110100",
       "00110011",
       "00110000",
       "00110000",
       "00110011",
       "00110100",
       "00111101",
       "01000011",
       "01001101",
       "01001100",
       "01010000",
       "01000011",
       "00111010",
       "00110100",
       "00100111",
       "00011100",
       "00110101",
       "00111011",
       "01001000",
       "01001110",
       "01001011",
       "01010011",
       "01010100",
       "01010101",
       "01010101",
       "01010110",
       "01010010",
       "01000101",
       "00111001",
       "00110110",
       "00110011",
       "00101101",
       "00100011",
       "00100110",
       "00100010",
       "00100000",
       "00011010",
       "00010110",
       "00010110",
       "00001010",
       "00011000",
       "00011101",
       "00010001",
       "00010111",
       "00010000",
       "00001111",
       "00011001",
       "00010001",
       "00010011",
       "00011110",
       "00110110",
       "00111011",
       "01001100",
       "01010010",
       "01010101",
       "01010100",
       "01011011",
       "01010111",
       "01010010",
       "01001110",
       "01000000",
       "00111000",
       "00110010",
       "00010001",
       "00011101",
       "00111100",
       "00111011",
       "01000010",
       "01001101",
       "01010110",
       "01000000",
       "00110110",
       "00110000",
       "00011101",
       "00100010",
       "00101001",
       "00011100",
       "00010000",
       "00001100",
       "00010001",
       "00010001",
       "00001111",
       "00001000",
       "00001111",
       "00010010",
       "00010111",
       "00100111",
       "00111010",
       "01000000",
       "00101101",
       "00111001",
       "00111110",
       "00110001",
       "00100110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00100011",
       "00010101",
       "00100110",
       "00111000",
       "00110011",
       "00110100",
       "00110001",
       "00110010",
       "00110010",
       "00110000",
       "00110001",
       "00110101",
       "00111010",
       "01000001",
       "01001100",
       "01001110",
       "01010010",
       "01001010",
       "01000000",
       "00111001",
       "00111011",
       "00100011",
       "00110011",
       "00111101",
       "01000111",
       "01010010",
       "01001101",
       "01010101",
       "01010100",
       "01010110",
       "01010111",
       "01010001",
       "01001111",
       "01000101",
       "00111010",
       "00111000",
       "00110011",
       "00101110",
       "00100011",
       "00100001",
       "00011011",
       "00010011",
       "00001101",
       "00001100",
       "00001101",
       "00001110",
       "00001011",
       "00001100",
       "00010010",
       "00010000",
       "00010010",
       "00010001",
       "00011000",
       "00001011",
       "00011001",
       "00011001",
       "00110000",
       "00111001",
       "01000101",
       "01010100",
       "01010101",
       "01011010",
       "01011000",
       "01010110",
       "01010100",
       "01001111",
       "00111111",
       "00111010",
       "00101000",
       "00010001",
       "00111001",
       "00111010",
       "01000001",
       "01001101",
       "01010010",
       "01010011",
       "01000011",
       "00110111",
       "00101111",
       "00101111",
       "00110110",
       "00111000",
       "00111001",
       "00101100",
       "00100000",
       "00001100",
       "00001100",
       "00010000",
       "00010001",
       "00001101",
       "00001010",
       "00010011",
       "00010100",
       "00100111",
       "01001101",
       "01000100",
       "00111001",
       "01000010",
       "00110111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001011",
       "00010001",
       "00101011",
       "00110111",
       "00110100",
       "00110111",
       "00110010",
       "00110110",
       "00110001",
       "00110001",
       "00110010",
       "00110011",
       "00111001",
       "01000010",
       "01001011",
       "01010001",
       "01010000",
       "01001111",
       "01001110",
       "01000000",
       "00111100",
       "00110110",
       "00111001",
       "00111110",
       "01001011",
       "01010001",
       "01001000",
       "01011001",
       "01011000",
       "01011001",
       "01010111",
       "01010101",
       "01010011",
       "01000111",
       "00111000",
       "00110110",
       "00110000",
       "00101111",
       "00100010",
       "00011100",
       "00010010",
       "00001100",
       "00001101",
       "00001010",
       "00001110",
       "00010000",
       "00001100",
       "00010100",
       "00001111",
       "00001100",
       "00010010",
       "00001101",
       "00010101",
       "00001011",
       "00010100",
       "00010111",
       "00101000",
       "00110101",
       "01000001",
       "01010011",
       "01010011",
       "01011011",
       "01010001",
       "01011000",
       "01010100",
       "01010011",
       "01000010",
       "00111111",
       "00100010",
       "00100011",
       "01000011",
       "00111111",
       "01001010",
       "01010011",
       "01011000",
       "01010010",
       "01000101",
       "00111000",
       "00110111",
       "00111000",
       "00110110",
       "00110011",
       "00110110",
       "00110100",
       "00110111",
       "00100011",
       "00010111",
       "00100000",
       "00100011",
       "00010000",
       "00000111",
       "00001101",
       "00010110",
       "00010111",
       "01000100",
       "01010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001101",
       "00010011",
       "00100110",
       "00110011",
       "00110110",
       "00110011",
       "00110101",
       "00110101",
       "00110100",
       "00110010",
       "00111001",
       "00110101",
       "00111010",
       "01000011",
       "01001100",
       "01010000",
       "01010000",
       "01010010",
       "01010100",
       "01001101",
       "01001000",
       "01000001",
       "00111110",
       "01000101",
       "01010110",
       "01010010",
       "01001011",
       "01011001",
       "01011000",
       "01011001",
       "01010111",
       "01010101",
       "01010001",
       "01000101",
       "00110111",
       "00110100",
       "00110011",
       "00101010",
       "00011110",
       "00011001",
       "00001101",
       "00001100",
       "00001110",
       "00001010",
       "00010000",
       "00001101",
       "00001101",
       "00010101",
       "00010000",
       "00001110",
       "00010110",
       "00001111",
       "00010011",
       "00001111",
       "00010000",
       "00011011",
       "00101010",
       "00110110",
       "00111111",
       "01010010",
       "01010100",
       "01010111",
       "01010110",
       "01011011",
       "01011001",
       "01011011",
       "01001010",
       "01000000",
       "00101101",
       "00110011",
       "01000001",
       "01000110",
       "01010010",
       "01010111",
       "01010110",
       "01010001",
       "01000010",
       "00111010",
       "00111001",
       "00111001",
       "00111001",
       "00111010",
       "00111000",
       "00110110",
       "00110101",
       "00110011",
       "00101100",
       "00110100",
       "00101101",
       "00011000",
       "00000110",
       "00010011",
       "00001100",
       "00011000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010001",
       "00010100",
       "00100101",
       "00110010",
       "00110110",
       "00110101",
       "00110011",
       "00110110",
       "00110101",
       "00110110",
       "00111010",
       "00111011",
       "01000010",
       "01000110",
       "01001110",
       "01010000",
       "01010011",
       "01010110",
       "01010101",
       "01011000",
       "01010100",
       "01010100",
       "01001101",
       "01010100",
       "01010111",
       "01010010",
       "01010010",
       "01011011",
       "01010110",
       "01011011",
       "01010110",
       "01010100",
       "01001111",
       "00111111",
       "00110110",
       "00110110",
       "00110011",
       "00100110",
       "00010101",
       "00010110",
       "00010010",
       "00001010",
       "00010000",
       "00001100",
       "00010010",
       "00001111",
       "00010001",
       "00010001",
       "00010100",
       "00010100",
       "00010010",
       "00010010",
       "00010100",
       "00010011",
       "00100000",
       "00011101",
       "00101111",
       "00111001",
       "01000001",
       "01001110",
       "01010111",
       "01010101",
       "01010111",
       "01011001",
       "01011101",
       "01011011",
       "01010100",
       "01000011",
       "00111100",
       "00111100",
       "01000101",
       "01010000",
       "01010100",
       "01010111",
       "01011100",
       "01001100",
       "01000100",
       "00111111",
       "00111010",
       "00111101",
       "01000100",
       "01000110",
       "01000101",
       "00111011",
       "00110111",
       "00110001",
       "00110100",
       "00110111",
       "00110111",
       "00100101",
       "00001011",
       "00001110",
       "00010000",
       "00001100",
       "00010101",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001101",
       "00010101",
       "00011110",
       "00110000",
       "00110010",
       "00110100",
       "00110000",
       "00111011",
       "00111011",
       "00111101",
       "01000000",
       "01001001",
       "01001000",
       "01001100",
       "01010101",
       "01010010",
       "01010010",
       "01010110",
       "01011001",
       "01011011",
       "01010100",
       "01011110",
       "01011110",
       "01011010",
       "01010101",
       "01010100",
       "01011000",
       "01011100",
       "01011101",
       "01011101",
       "01011001",
       "01011000",
       "01001110",
       "00111000",
       "00110101",
       "00110100",
       "00110010",
       "00110011",
       "00101110",
       "00101001",
       "00011011",
       "00001100",
       "00001110",
       "00001101",
       "00010001",
       "00010011",
       "00010010",
       "00010100",
       "00010111",
       "00011100",
       "00010110",
       "00011010",
       "00010011",
       "00010111",
       "00011111",
       "00100000",
       "00101111",
       "00111000",
       "00111100",
       "01001001",
       "01010100",
       "01011001",
       "01010111",
       "01011100",
       "01011101",
       "01011110",
       "01011101",
       "01001101",
       "01000111",
       "01000110",
       "01010011",
       "01011001",
       "01011011",
       "01011010",
       "01010111",
       "01001000",
       "01001101",
       "01001010",
       "01000101",
       "01000110",
       "01001000",
       "01001010",
       "01001001",
       "01000001",
       "00111110",
       "00111001",
       "00111010",
       "00110011",
       "00111010",
       "00101000",
       "00001100",
       "00001010",
       "00010001",
       "00001110",
       "00011001",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001011",
       "00001111",
       "00011010",
       "00101000",
       "00110101",
       "00110001",
       "00110101",
       "00111110",
       "01000011",
       "01000111",
       "01001101",
       "01001111",
       "01001101",
       "01010000",
       "01010101",
       "01010101",
       "01010110",
       "01011001",
       "01011011",
       "01011011",
       "01011000",
       "01010111",
       "01011010",
       "01011101",
       "01011011",
       "01010111",
       "01011100",
       "01011100",
       "01011010",
       "01011010",
       "01011011",
       "01011010",
       "01001011",
       "00111001",
       "00110101",
       "00110011",
       "00111000",
       "00110111",
       "00111110",
       "00111010",
       "00101010",
       "00010011",
       "00010011",
       "00011110",
       "00011001",
       "00010110",
       "00001010",
       "00011100",
       "00110001",
       "00110110",
       "00111010",
       "00111001",
       "00101001",
       "00100000",
       "00100100",
       "00110000",
       "00110010",
       "00111011",
       "00110111",
       "01001110",
       "01010110",
       "01011011",
       "01011011",
       "01100000",
       "01011011",
       "01100001",
       "01011010",
       "01010101",
       "01010111",
       "01011011",
       "01011001",
       "01011010",
       "01011001",
       "01011101",
       "01001110",
       "01001100",
       "01010100",
       "01001101",
       "01001100",
       "01010001",
       "01001101",
       "01010000",
       "01001110",
       "01001011",
       "01000111",
       "01000010",
       "00111100",
       "00110111",
       "00110101",
       "00101001",
       "00001011",
       "00001110",
       "00001100",
       "00010011",
       "00010011",
       "00010111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001011",
       "00001000",
       "00001011",
       "00010001",
       "00011110",
       "00101111",
       "00110111",
       "00110111",
       "00111001",
       "00111101",
       "01000101",
       "01000111",
       "01010000",
       "01001101",
       "01010000",
       "01010001",
       "01010110",
       "01010111",
       "01011001",
       "01010101",
       "01011100",
       "01011010",
       "01011011",
       "01010111",
       "01011111",
       "01011110",
       "01011011",
       "01011011",
       "01011010",
       "01010010",
       "01011001",
       "01011000",
       "01011010",
       "01001110",
       "01000010",
       "00111001",
       "00110111",
       "00111001",
       "00110110",
       "00110110",
       "00111100",
       "00111101",
       "00101000",
       "00010111",
       "00101101",
       "00100110",
       "00010010",
       "00010000",
       "00110001",
       "00111110",
       "00111111",
       "01000010",
       "01000000",
       "00111110",
       "00111000",
       "00110110",
       "00110100",
       "00111001",
       "00111100",
       "00111101",
       "01010101",
       "01011010",
       "01011010",
       "01011100",
       "01011101",
       "01011100",
       "01011101",
       "01011001",
       "01001110",
       "01011101",
       "01011011",
       "01011001",
       "01010110",
       "01011100",
       "01011000",
       "01001110",
       "01010100",
       "01010110",
       "01010010",
       "01010100",
       "01010110",
       "01010001",
       "01001110",
       "01010010",
       "01001001",
       "01001101",
       "01000011",
       "00111101",
       "00111000",
       "00111001",
       "00011111",
       "00001101",
       "00010010",
       "00001111",
       "00010001",
       "00001101",
       "00010111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001110",
       "00001111",
       "00001100",
       "00001100",
       "00001001",
       "00001111",
       "00011101",
       "00110010",
       "00110101",
       "00111010",
       "00110101",
       "00110111",
       "00110101",
       "00111111",
       "01000101",
       "01010011",
       "01010011",
       "01010111",
       "01010110",
       "01011000",
       "01010111",
       "01011100",
       "01011101",
       "01011110",
       "01011011",
       "01011100",
       "01011111",
       "01011101",
       "01011110",
       "01010111",
       "01011001",
       "01011001",
       "01010110",
       "01011010",
       "01010011",
       "01001110",
       "01000100",
       "01000100",
       "01000101",
       "01000110",
       "00111110",
       "00111110",
       "00111110",
       "00111001",
       "00101001",
       "00101110",
       "00110111",
       "00100010",
       "00010111",
       "00111011",
       "00110100",
       "00111111",
       "01000000",
       "00111000",
       "00111001",
       "00111010",
       "00111100",
       "00111001",
       "00111111",
       "01000010",
       "01001011",
       "01010111",
       "01011011",
       "01011001",
       "01011010",
       "01011111",
       "01011101",
       "01011111",
       "01010011",
       "01001010",
       "01011111",
       "01010111",
       "01011101",
       "01011001",
       "01011110",
       "01010110",
       "01011001",
       "01010110",
       "01011001",
       "01010101",
       "01010010",
       "01010001",
       "01010010",
       "01001111",
       "01010011",
       "01001100",
       "01001010",
       "00111110",
       "00111100",
       "00110111",
       "00110110",
       "00010101",
       "00001110",
       "00010010",
       "00010010",
       "00010100",
       "00010101",
       "00010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010001",
       "00010001",
       "00010001",
       "00010010",
       "00001111",
       "00001100",
       "00001010",
       "00001101",
       "00010110",
       "00100001",
       "00100111",
       "00101110",
       "00110011",
       "00110111",
       "00110111",
       "00111011",
       "01000000",
       "01001111",
       "01010111",
       "01011011",
       "01011010",
       "01011100",
       "01011011",
       "01100000",
       "01011110",
       "01011101",
       "01011100",
       "01011111",
       "01011011",
       "01011101",
       "01011010",
       "01011110",
       "01011100",
       "01011110",
       "01010111",
       "01001111",
       "01011010",
       "01011001",
       "01010101",
       "01010100",
       "01010001",
       "01000110",
       "00111101",
       "00111010",
       "00111010",
       "00111100",
       "00111000",
       "00111111",
       "00110101",
       "00011100",
       "00111000",
       "00111001",
       "01000101",
       "01001111",
       "01000100",
       "00111110",
       "00111011",
       "01000011",
       "01000101",
       "01001100",
       "01010100",
       "01010111",
       "01011000",
       "01011110",
       "01011100",
       "01011100",
       "01011110",
       "01011110",
       "01100001",
       "01001110",
       "01001111",
       "01011111",
       "01011110",
       "01011111",
       "01011101",
       "01011010",
       "01011010",
       "01011111",
       "01011010",
       "01011000",
       "01010011",
       "01010000",
       "01010001",
       "01010010",
       "01010001",
       "01010001",
       "01001011",
       "01000101",
       "00111110",
       "00111010",
       "00111001",
       "00100010",
       "00010000",
       "00010100",
       "00001111",
       "00011011",
       "00011111",
       "00101010",
       "00011110",
       "00010111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00011000",
       "00001101",
       "00010101",
       "00001010",
       "00001111",
       "00001011",
       "00010001",
       "00010001",
       "00011101",
       "00011110",
       "00100100",
       "00100101",
       "00100100",
       "00011111",
       "00101010",
       "00110100",
       "00111010",
       "00110111",
       "01000100",
       "01001110",
       "01010100",
       "01011000",
       "01011100",
       "01011010",
       "01100000",
       "01011100",
       "01011101",
       "01011001",
       "01011111",
       "01011111",
       "01011101",
       "01011101",
       "01100000",
       "01100000",
       "01011101",
       "01010101",
       "01010000",
       "01011000",
       "01011111",
       "01011101",
       "01011001",
       "01011100",
       "01010110",
       "01001011",
       "00111111",
       "00111111",
       "00111101",
       "00111111",
       "00111100",
       "00111011",
       "00100100",
       "00110111",
       "00111110",
       "01000110",
       "01010010",
       "01010001",
       "01001100",
       "01001011",
       "01010010",
       "01011001",
       "01100000",
       "01100000",
       "01011100",
       "01011010",
       "01100000",
       "01100010",
       "01100001",
       "01011100",
       "01011110",
       "01011101",
       "01010111",
       "01011001",
       "01011110",
       "01100001",
       "01011111",
       "01010110",
       "01011111",
       "01011101",
       "01100000",
       "01011011",
       "01011001",
       "01010110",
       "01010100",
       "01010110",
       "01010010",
       "01001010",
       "01001010",
       "01000001",
       "00111010",
       "00111011",
       "00111000",
       "00101110",
       "00010101",
       "00001110",
       "00001110",
       "00011110",
       "00100100",
       "00101111",
       "00110101",
       "00110101",
       "00101011",
       "00011110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010111",
       "00010001",
       "00010000",
       "00010110",
       "00001111",
       "00001011",
       "00010001",
       "00011000",
       "00100101",
       "00110010",
       "00110101",
       "00110101",
       "00110110",
       "00110011",
       "00101010",
       "00011101",
       "00011011",
       "00100111",
       "00111000",
       "00111000",
       "01000011",
       "01001111",
       "01010111",
       "01011000",
       "01011101",
       "01011110",
       "01011111",
       "01011110",
       "01100000",
       "01011110",
       "01011111",
       "01011101",
       "01011111",
       "01011101",
       "01011101",
       "01011111",
       "01011101",
       "01010011",
       "01010100",
       "01011100",
       "01011101",
       "01011101",
       "01011101",
       "01011101",
       "01011100",
       "01010101",
       "01010110",
       "01001110",
       "01000101",
       "01000001",
       "01000000",
       "00011111",
       "00101110",
       "01000000",
       "01000011",
       "01010110",
       "01011011",
       "01011010",
       "01010101",
       "01010110",
       "01011101",
       "01100010",
       "01100001",
       "01011111",
       "01011110",
       "01011111",
       "01100001",
       "01100001",
       "01011111",
       "01011111",
       "01011100",
       "01011010",
       "01011100",
       "01100100",
       "01100000",
       "01011000",
       "01011011",
       "01100000",
       "01011000",
       "01011100",
       "01011001",
       "01011000",
       "01010001",
       "01001101",
       "01000110",
       "01000011",
       "00111011",
       "00111001",
       "00111000",
       "00111000",
       "00111011",
       "00110101",
       "00011100",
       "00010011",
       "00011001",
       "00011010",
       "00101101",
       "00110001",
       "00111010",
       "00111010",
       "01000000",
       "00110101",
       "00110100",
       "00010101",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001000",
       "00010110",
       "01000000",
       "00110001",
       "00101110",
       "00110011",
       "01010010",
       "00110010",
       "00010001",
       "00010011",
       "00010100",
       "00010110",
       "00011101",
       "00011101",
       "00011101",
       "00011100",
       "00101001",
       "00110100",
       "00110100",
       "00110101",
       "00110000",
       "00110011",
       "00110110",
       "00111010",
       "00110101",
       "00101110",
       "00011011",
       "00100011",
       "00110001",
       "00111110",
       "01010001",
       "01011010",
       "01011010",
       "01011101",
       "01011111",
       "01100011",
       "01011100",
       "01100010",
       "01100000",
       "01011111",
       "01011110",
       "01100000",
       "01011010",
       "01011101",
       "01011011",
       "01010101",
       "01010010",
       "01011000",
       "01011101",
       "01011010",
       "01011001",
       "01010111",
       "01100001",
       "01100011",
       "01100100",
       "01011100",
       "01010011",
       "01000101",
       "00111101",
       "00111010",
       "00011101",
       "00110011",
       "00111110",
       "01000111",
       "01011000",
       "01100010",
       "01100101",
       "01011111",
       "01011100",
       "01011100",
       "01011011",
       "01011111",
       "01100001",
       "01011101",
       "01011101",
       "01011100",
       "01100010",
       "01100011",
       "01011111",
       "01011110",
       "01011001",
       "01011101",
       "01011111",
       "01011010",
       "01011001",
       "01011101",
       "01100000",
       "01011011",
       "01011010",
       "01010100",
       "01001111",
       "01000101",
       "00111101",
       "00111001",
       "00111000",
       "00110101",
       "00111000",
       "00111010",
       "00111110",
       "00110000",
       "00100000",
       "00010100",
       "00011100",
       "00101001",
       "00110010",
       "00110110",
       "00111100",
       "00111011",
       "00111111",
       "00111100",
       "00111100",
       "00110111",
       "00110011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001000",
       "00101110",
       "00110111",
       "00101100",
       "00101011",
       "01001001",
       "01000011",
       "00010100",
       "00010011",
       "00011100",
       "00100101",
       "00101001",
       "00101110",
       "00101110",
       "00110010",
       "00110000",
       "00110110",
       "00110111",
       "00111001",
       "00110111",
       "00111011",
       "00111011",
       "00111000",
       "00110010",
       "00110101",
       "00111001",
       "00110111",
       "00101100",
       "00110110",
       "00111101",
       "01001100",
       "01010110",
       "01011110",
       "01011011",
       "01011101",
       "01011110",
       "01011101",
       "01011111",
       "01100000",
       "01011110",
       "01100000",
       "01011110",
       "01011110",
       "01011101",
       "01010110",
       "01001101",
       "01001101",
       "01011000",
       "01011111",
       "01100000",
       "01011111",
       "01100000",
       "01101000",
       "01011111",
       "01011111",
       "01011000",
       "01001111",
       "00111100",
       "01000000",
       "00110110",
       "00100101",
       "01000000",
       "00111111",
       "01010001",
       "01011001",
       "01100011",
       "01100101",
       "01101001",
       "01100100",
       "01100101",
       "01100010",
       "01011100",
       "01100000",
       "01011010",
       "01011010",
       "01011101",
       "01100000",
       "01100100",
       "01100000",
       "01011011",
       "01011110",
       "01100000",
       "01011100",
       "01011010",
       "01011111",
       "01011010",
       "01100010",
       "01011001",
       "01010100",
       "01001001",
       "01000011",
       "00111101",
       "00111011",
       "00111001",
       "00111010",
       "00111010",
       "00111011",
       "00110000",
       "00101001",
       "00011000",
       "00011011",
       "00011101",
       "00101100",
       "00110010",
       "00111001",
       "00111000",
       "00111111",
       "00111010",
       "00111111",
       "00111101",
       "01000010",
       "00111001",
       "00111011",
       "00001100",
       "00101110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001001",
       "00110111",
       "00110010",
       "00101100",
       "00100111",
       "00111110",
       "00100010",
       "00010000",
       "00100010",
       "00101010",
       "00111001",
       "00110111",
       "00111010",
       "00111001",
       "00110111",
       "00111001",
       "00111101",
       "00111001",
       "00111011",
       "00111110",
       "01000111",
       "01001010",
       "01001101",
       "01000110",
       "00111100",
       "00110010",
       "00111000",
       "00111010",
       "00111101",
       "01000100",
       "01010100",
       "01011001",
       "01100010",
       "01100010",
       "01100000",
       "01011111",
       "01011111",
       "01011101",
       "01100011",
       "01100000",
       "01100000",
       "01011100",
       "01100101",
       "01011111",
       "01011100",
       "01010001",
       "01001111",
       "01010111",
       "01011110",
       "01100000",
       "01100101",
       "01100001",
       "01100011",
       "01100001",
       "01100011",
       "01100001",
       "01011011",
       "01000001",
       "01000001",
       "00101011",
       "00101011",
       "01000000",
       "01000001",
       "01010110",
       "01100000",
       "01100010",
       "01101000",
       "01101000",
       "01100100",
       "01100010",
       "01100101",
       "01011110",
       "01100000",
       "01011111",
       "01011010",
       "01100010",
       "01011111",
       "01011110",
       "01011011",
       "01011110",
       "01100000",
       "01011111",
       "01100001",
       "01011111",
       "01100010",
       "01100010",
       "01100000",
       "01010101",
       "01001010",
       "01000001",
       "01000000",
       "00111110",
       "00111101",
       "00111010",
       "00110000",
       "00100110",
       "00100110",
       "00011001",
       "00010110",
       "00011011",
       "00100110",
       "00101110",
       "00111010",
       "00111010",
       "00111110",
       "00111101",
       "00111111",
       "00111001",
       "00111101",
       "00111111",
       "01000010",
       "01000000",
       "00111011",
       "00011000",
       "00010001",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00011001",
       "00111011",
       "00110001",
       "00110001",
       "00101110",
       "00101010",
       "00010111",
       "00100100",
       "00110000",
       "00110111",
       "00111010",
       "00111010",
       "00111001",
       "00111000",
       "00111000",
       "00111001",
       "00111101",
       "00111111",
       "01000011",
       "01000111",
       "01001101",
       "01001111",
       "01010110",
       "01010101",
       "01001110",
       "01000111",
       "01000101",
       "01000100",
       "01001011",
       "01010110",
       "01100001",
       "01011101",
       "01011100",
       "01011010",
       "01011111",
       "01011111",
       "01100000",
       "01100000",
       "01100001",
       "01100001",
       "01100100",
       "01100011",
       "01100011",
       "01011110",
       "01011110",
       "01011001",
       "01011001",
       "01011010",
       "01011100",
       "01011111",
       "01100010",
       "01011101",
       "01100011",
       "01010110",
       "01010010",
       "01010011",
       "01010110",
       "01000101",
       "01000010",
       "00101011",
       "00110000",
       "01000001",
       "01000000",
       "01011100",
       "01011110",
       "01011110",
       "01101010",
       "01101011",
       "01100110",
       "01100011",
       "01011111",
       "01100000",
       "01100000",
       "01100101",
       "01011100",
       "01100010",
       "01100001",
       "01011101",
       "01011110",
       "01100101",
       "01100000",
       "01100001",
       "01011110",
       "01011011",
       "01100001",
       "01100110",
       "01100000",
       "01011000",
       "01000011",
       "00111110",
       "00111100",
       "00111101",
       "00110111",
       "00110101",
       "00100100",
       "00010111",
       "00010100",
       "00011001",
       "00011111",
       "00101001",
       "00101110",
       "00111100",
       "00111101",
       "00111100",
       "00111011",
       "00111111",
       "00111101",
       "00111100",
       "00111110",
       "01000000",
       "00111101",
       "01000000",
       "00111010",
       "00100110",
       "00000101",
       "00110011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001100",
       "00101000",
       "00111001",
       "00110100",
       "00110101",
       "00101011",
       "00011101",
       "00100111",
       "00110100",
       "00110111",
       "00111101",
       "00111011",
       "00111101",
       "01000000",
       "01000010",
       "01000100",
       "01000101",
       "01000011",
       "01000110",
       "01001101",
       "01010000",
       "01001111",
       "01010000",
       "01010110",
       "01010110",
       "01010111",
       "01010111",
       "01011011",
       "01011001",
       "01011010",
       "01011100",
       "01011100",
       "01011001",
       "01010110",
       "01010011",
       "01010101",
       "01011000",
       "01100000",
       "01100001",
       "01100000",
       "01100011",
       "01100000",
       "01100101",
       "01100100",
       "01100001",
       "01100100",
       "01011101",
       "01011011",
       "01011111",
       "01100001",
       "01100010",
       "01011110",
       "01100010",
       "01011011",
       "01000101",
       "01000001",
       "01000101",
       "01000010",
       "00111111",
       "00111110",
       "00011111",
       "00011011",
       "00111011",
       "00111101",
       "01001101",
       "01010011",
       "01011000",
       "01100110",
       "01101001",
       "01100111",
       "01100011",
       "01011111",
       "01011101",
       "01100000",
       "01100001",
       "01100001",
       "01100100",
       "01100001",
       "01100000",
       "01100011",
       "01100010",
       "01100001",
       "01100011",
       "01011111",
       "01011101",
       "01100010",
       "01100100",
       "01100001",
       "01011010",
       "01000101",
       "00111100",
       "00110111",
       "00111001",
       "00110100",
       "00110010",
       "00100101",
       "00010100",
       "00001110",
       "00011110",
       "00100100",
       "00101111",
       "00110100",
       "00111010",
       "00111001",
       "00111010",
       "00111100",
       "01000001",
       "00111010",
       "01000000",
       "00111111",
       "01000011",
       "00111110",
       "01000001",
       "00111011",
       "00111010",
       "00001101",
       "00010100",
       "01000010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010110",
       "00100100",
       "00101111",
       "00110000",
       "00101011",
       "00100101",
       "00100101",
       "00110110",
       "00111110",
       "00111011",
       "00111110",
       "01000011",
       "01000110",
       "01001101",
       "01010000",
       "01010000",
       "01001110",
       "01010011",
       "01010000",
       "01010000",
       "01010001",
       "01010101",
       "01010100",
       "01010100",
       "01010111",
       "01010111",
       "01011010",
       "01011010",
       "01011001",
       "01011011",
       "01100000",
       "01011100",
       "01100001",
       "01011111",
       "01100010",
       "01011101",
       "01100000",
       "01100000",
       "01100001",
       "01100001",
       "01100011",
       "01100000",
       "01100101",
       "01100001",
       "01100001",
       "01100010",
       "01100001",
       "01011011",
       "01011101",
       "01011111",
       "01100010",
       "01011110",
       "01100010",
       "01010110",
       "01000110",
       "00111001",
       "01000000",
       "00111011",
       "01000011",
       "00101111",
       "00101101",
       "00011111",
       "00101000",
       "01001001",
       "00111101",
       "01000011",
       "01000111",
       "01011111",
       "01100100",
       "01101000",
       "01100100",
       "01100100",
       "01011111",
       "01011111",
       "01100010",
       "01100010",
       "01100010",
       "01100001",
       "01011101",
       "01100001",
       "01100010",
       "01100011",
       "01100010",
       "01100010",
       "01100100",
       "01100100",
       "01100010",
       "01100010",
       "01011001",
       "01001000",
       "01000001",
       "00111011",
       "00101111",
       "00101000",
       "00100101",
       "00100000",
       "00010100",
       "00010100",
       "00011110",
       "00100101",
       "00110000",
       "00111000",
       "00111010",
       "00111011",
       "00111100",
       "01000001",
       "00111101",
       "00111100",
       "01000000",
       "01000010",
       "01001000",
       "01000110",
       "00111111",
       "01000001",
       "00111100",
       "00110001",
       "00000110",
       "00111000",
       "00101111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010001",
       "00101001",
       "00101000",
       "00110001",
       "00010111",
       "00100110",
       "00110110",
       "00111110",
       "01000001",
       "00111101",
       "01000100",
       "01001110",
       "01010110",
       "01010111",
       "01011001",
       "01010101",
       "01010011",
       "01010110",
       "01010110",
       "01010100",
       "01010010",
       "01010011",
       "01010011",
       "01010100",
       "01010000",
       "01010000",
       "01011001",
       "01010111",
       "01011010",
       "01011110",
       "01100001",
       "01011101",
       "01100000",
       "01100000",
       "01100100",
       "01100011",
       "01100010",
       "01011111",
       "01100001",
       "01100011",
       "01100010",
       "01100010",
       "01100001",
       "01011111",
       "01011111",
       "01100011",
       "01100001",
       "01011011",
       "01011110",
       "01011100",
       "01100100",
       "01100001",
       "01100101",
       "01100001",
       "01011101",
       "01000010",
       "00110111",
       "00100101",
       "00110010",
       "00100010",
       "00110010",
       "00101010",
       "00001011",
       "00111001",
       "00110110",
       "01001011",
       "01010011",
       "01100011",
       "01100100",
       "01100111",
       "01100101",
       "01100101",
       "01100010",
       "01011110",
       "01100011",
       "01011110",
       "01011101",
       "01100010",
       "01100000",
       "01100000",
       "01100010",
       "01100100",
       "01100010",
       "01011110",
       "01100000",
       "01011110",
       "01100001",
       "01100101",
       "01100000",
       "01010011",
       "01000110",
       "01000011",
       "00111011",
       "00110000",
       "00100001",
       "00010010",
       "00010001",
       "00011001",
       "00010110",
       "00100000",
       "00101010",
       "00110110",
       "00111100",
       "01000010",
       "00111111",
       "01000000",
       "00111001",
       "00111110",
       "01000010",
       "01000110",
       "01001100",
       "01001110",
       "01000000",
       "01000011",
       "00111001",
       "01000001",
       "00010011",
       "00011110",
       "00111100",
       "00100100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010001",
       "00101101",
       "00101101",
       "00110110",
       "00010001",
       "00101011",
       "00111101",
       "01000010",
       "01000010",
       "01000111",
       "01010001",
       "01010110",
       "01011000",
       "01010010",
       "01010001",
       "01010001",
       "01010010",
       "01010010",
       "01010010",
       "01010110",
       "01010111",
       "01001100",
       "01000011",
       "01000010",
       "01000111",
       "01001111",
       "01010010",
       "01010111",
       "01011110",
       "01100000",
       "01011101",
       "01011111",
       "01011101",
       "01011111",
       "01011101",
       "01011111",
       "01011110",
       "01100001",
       "01100000",
       "01100001",
       "01100000",
       "01100100",
       "01100000",
       "01011111",
       "01011100",
       "01011101",
       "01011101",
       "01011110",
       "01011111",
       "01100000",
       "01100110",
       "01100101",
       "01100010",
       "01100101",
       "01101000",
       "01101010",
       "01100100",
       "01001101",
       "01001000",
       "01000101",
       "00111110",
       "01000100",
       "01000100",
       "01000101",
       "01011000",
       "01101000",
       "01101011",
       "01100110",
       "01100010",
       "01100111",
       "01100110",
       "01100100",
       "01100001",
       "01100011",
       "01100010",
       "01011101",
       "01011101",
       "01011011",
       "01011101",
       "01100100",
       "01100010",
       "01100100",
       "01100001",
       "01011011",
       "01011101",
       "01011100",
       "01100100",
       "01100100",
       "01100100",
       "01100010",
       "01010110",
       "01000110",
       "01000111",
       "01000001",
       "00111010",
       "00101111",
       "00100101",
       "00100100",
       "00101001",
       "00101000",
       "00101011",
       "00101011",
       "00101111",
       "00111010",
       "00111111",
       "00111111",
       "00111111",
       "01000000",
       "01001001",
       "01001101",
       "01001111",
       "01010100",
       "01001001",
       "01000011",
       "00111101",
       "00111110",
       "00110001",
       "00001011",
       "00110111",
       "00011101",
       "00100100",
       "00101100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00100100",
       "00110101",
       "00111000",
       "00001110",
       "00110011",
       "00111111",
       "01000010",
       "01000100",
       "01010100",
       "01010110",
       "01010110",
       "01010000",
       "01000101",
       "01000001",
       "01000010",
       "01001000",
       "01010000",
       "01001111",
       "01001111",
       "01001111",
       "01000111",
       "00111110",
       "00111110",
       "01000100",
       "01001100",
       "01010101",
       "01011110",
       "01011010",
       "01011110",
       "01011110",
       "01011101",
       "01011101",
       "01100010",
       "01011110",
       "01100010",
       "01100101",
       "01100011",
       "01100011",
       "01011111",
       "01100001",
       "01100100",
       "01100001",
       "01010101",
       "01010111",
       "01011010",
       "01011010",
       "01011110",
       "01011000",
       "01011011",
       "01011101",
       "01100101",
       "01100101",
       "01101001",
       "01100110",
       "01100111",
       "01101110",
       "01111000",
       "01110110",
       "01110101",
       "01110001",
       "01110101",
       "01111110",
       "01110101",
       "01101101",
       "01100110",
       "01101010",
       "01101000",
       "01101010",
       "01100011",
       "01100110",
       "01100001",
       "01100001",
       "01011000",
       "01010110",
       "01010011",
       "01010111",
       "01001100",
       "01011001",
       "01100010",
       "01100000",
       "01100000",
       "01100010",
       "01100001",
       "01100000",
       "01100010",
       "01100101",
       "01100110",
       "01100100",
       "01100001",
       "01100001",
       "01010110",
       "01001111",
       "01000110",
       "01000011",
       "01000101",
       "01000010",
       "00111001",
       "00111110",
       "00111010",
       "00110100",
       "00101101",
       "00100110",
       "00101011",
       "00111001",
       "00111111",
       "01000011",
       "00111111",
       "01001100",
       "01010010",
       "01011001",
       "01011000",
       "01010100",
       "01000110",
       "01000000",
       "00111110",
       "01000001",
       "00011000",
       "00100110",
       "00011010",
       "00110000",
       "00101101",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00101110",
       "00101001",
       "00001100",
       "00110100",
       "01000001",
       "01000010",
       "01001000",
       "01010101",
       "01010111",
       "01010011",
       "01001001",
       "00111010",
       "00111000",
       "00111001",
       "00111110",
       "01001000",
       "01001001",
       "01001010",
       "01000101",
       "00111110",
       "01000010",
       "01000000",
       "01000101",
       "01010000",
       "01010111",
       "01011101",
       "01011110",
       "01011111",
       "01011101",
       "01011111",
       "01100010",
       "01100011",
       "01100010",
       "01100010",
       "01100110",
       "01100010",
       "01100011",
       "01100010",
       "01100000",
       "01100001",
       "01100111",
       "01011100",
       "01010101",
       "01010101",
       "01001110",
       "01000101",
       "01010100",
       "01011100",
       "01011100",
       "01100000",
       "01100100",
       "01100010",
       "01100101",
       "01100011",
       "01100110",
       "01101111",
       "01101001",
       "01101010",
       "01101101",
       "01101100",
       "01101101",
       "01101101",
       "01101000",
       "01101011",
       "01101110",
       "01101011",
       "01101011",
       "01101010",
       "01101010",
       "01011010",
       "01000110",
       "00110010",
       "00111010",
       "01010000",
       "01011000",
       "01010011",
       "01011011",
       "01100011",
       "01100001",
       "01100011",
       "01100011",
       "01100101",
       "01100100",
       "01100101",
       "01100101",
       "01100010",
       "01100011",
       "01100111",
       "01100011",
       "01100000",
       "01100000",
       "01011010",
       "01010001",
       "01001001",
       "01000111",
       "01000100",
       "01000001",
       "01000001",
       "01000000",
       "00111100",
       "00101010",
       "00100100",
       "00110101",
       "01000001",
       "01000100",
       "01000000",
       "01001011",
       "01010001",
       "01011100",
       "01011011",
       "01011000",
       "01001001",
       "01000011",
       "00111111",
       "01000001",
       "00110000",
       "00011011",
       "00011011",
       "00100110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00011010",
       "00001000",
       "00110111",
       "01000010",
       "01000111",
       "01001001",
       "01010011",
       "01010110",
       "01001110",
       "01000101",
       "00111111",
       "00110001",
       "00111001",
       "00111010",
       "00111101",
       "01000000",
       "01000010",
       "00111110",
       "00111101",
       "00111100",
       "00111001",
       "01000100",
       "01010011",
       "01011100",
       "01011110",
       "01100001",
       "01100000",
       "01100000",
       "01100110",
       "01100100",
       "01100010",
       "01011111",
       "01100000",
       "01100011",
       "01100011",
       "01100011",
       "01100001",
       "01011111",
       "01100100",
       "01101000",
       "01100010",
       "01010101",
       "01010010",
       "01001001",
       "00111010",
       "01000010",
       "01010001",
       "01011010",
       "01011000",
       "01100010",
       "01100011",
       "01101000",
       "01100110",
       "01100111",
       "01101001",
       "01101110",
       "01101111",
       "01101010",
       "01101100",
       "01110000",
       "01101100",
       "01100111",
       "01101100",
       "01101100",
       "01101111",
       "01101011",
       "01011110",
       "01000010",
       "00100110",
       "00010110",
       "00001111",
       "00101111",
       "01001011",
       "01010000",
       "01011110",
       "01011110",
       "01100110",
       "01100001",
       "01100010",
       "01100100",
       "01100010",
       "01100001",
       "01100001",
       "01100011",
       "01100010",
       "01100010",
       "01100110",
       "01100111",
       "01100100",
       "01100010",
       "01100010",
       "01100011",
       "01011100",
       "01011100",
       "01010111",
       "01010001",
       "01001101",
       "01000101",
       "01000010",
       "00110101",
       "00101000",
       "00101110",
       "01000000",
       "01000010",
       "01000001",
       "01001010",
       "01010100",
       "01010110",
       "01010111",
       "01010010",
       "01001101",
       "01000001",
       "01000010",
       "00111111",
       "01000000",
       "00011111",
       "00011110",
       "00001110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00100010",
       "00001000",
       "00110100",
       "00111101",
       "01001000",
       "01000111",
       "01010010",
       "01010100",
       "01001110",
       "01000010",
       "01000001",
       "00101100",
       "00110001",
       "00110111",
       "00111011",
       "00111110",
       "00111110",
       "00111101",
       "00111010",
       "00111011",
       "00111101",
       "01001011",
       "01011000",
       "01100000",
       "01011101",
       "01011110",
       "01100011",
       "01100001",
       "01100100",
       "01100011",
       "01100000",
       "01011100",
       "01100010",
       "01100011",
       "01100111",
       "01100100",
       "01100010",
       "01100010",
       "01100010",
       "01100110",
       "01010111",
       "01001110",
       "01010001",
       "01000101",
       "01000100",
       "00111101",
       "00101000",
       "00011111",
       "00101010",
       "00111100",
       "01010010",
       "01100100",
       "01101010",
       "01101110",
       "01101000",
       "01101100",
       "01101110",
       "01101100",
       "01101100",
       "01101000",
       "01101010",
       "01101011",
       "01101101",
       "01101011",
       "01010111",
       "00111011",
       "00100000",
       "00001100",
       "00000111",
       "00001001",
       "00001110",
       "00111010",
       "01001000",
       "01001000",
       "01010011",
       "01100011",
       "01100101",
       "01100011",
       "01100011",
       "01100100",
       "01100010",
       "01100001",
       "01100001",
       "01100000",
       "01100011",
       "01100110",
       "01100111",
       "01100100",
       "01101000",
       "01100101",
       "01100011",
       "01100000",
       "01100000",
       "01100011",
       "01100010",
       "01011100",
       "01010111",
       "01001100",
       "01000001",
       "01000000",
       "00110111",
       "00110011",
       "01000000",
       "01000101",
       "01001000",
       "01001100",
       "01011001",
       "01010110",
       "01011010",
       "01010011",
       "01010011",
       "01000110",
       "01000100",
       "00111011",
       "01000000",
       "00101101",
       "00011111",
       "00001000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00100101",
       "00001011",
       "00101011",
       "00111010",
       "01000100",
       "01000011",
       "01001111",
       "01011001",
       "01001111",
       "01000100",
       "01000000",
       "00110111",
       "00100111",
       "00101101",
       "00111001",
       "00111101",
       "00111011",
       "00111110",
       "00110111",
       "00111010",
       "01000011",
       "01010011",
       "01011000",
       "01011011",
       "01011100",
       "01011100",
       "01100000",
       "01011111",
       "01011100",
       "01011111",
       "01011110",
       "01100010",
       "01100100",
       "01100011",
       "01100011",
       "01100010",
       "01100100",
       "01100100",
       "01100001",
       "01100101",
       "01010111",
       "01001001",
       "01001001",
       "01000110",
       "01000100",
       "01001011",
       "00110011",
       "00001000",
       "00001010",
       "00000111",
       "00011010",
       "00100000",
       "00111010",
       "01010100",
       "01100111",
       "01110000",
       "01100111",
       "01100101",
       "01100110",
       "01101001",
       "01101110",
       "01011110",
       "01001011",
       "00110000",
       "00011001",
       "00001100",
       "00001110",
       "00010001",
       "00010001",
       "00010000",
       "00101111",
       "01001010",
       "01001100",
       "01001111",
       "01010100",
       "01100100",
       "01100101",
       "01100101",
       "01100101",
       "01100001",
       "01100010",
       "01100000",
       "01011101",
       "01011011",
       "01010111",
       "01100000",
       "01100101",
       "01100011",
       "01100110",
       "01100111",
       "01100111",
       "01100010",
       "01100011",
       "01100000",
       "01011111",
       "01011110",
       "01011001",
       "01011001",
       "01001101",
       "01000110",
       "01000010",
       "00111101",
       "01000101",
       "01000111",
       "01001011",
       "01010011",
       "01011011",
       "01011010",
       "01011101",
       "01011000",
       "01010101",
       "01001101",
       "01000010",
       "00111110",
       "00111110",
       "00111000",
       "00100000",
       "00010100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00100100",
       "00010100",
       "00101000",
       "00110001",
       "01000001",
       "01000010",
       "01001100",
       "01011001",
       "01010100",
       "01001010",
       "01000010",
       "00111101",
       "00101111",
       "00100010",
       "00110101",
       "00111101",
       "00111100",
       "00111111",
       "01000000",
       "00111101",
       "01000011",
       "01010001",
       "01010001",
       "01011011",
       "01011011",
       "01011110",
       "01011111",
       "01011111",
       "01011110",
       "01100011",
       "01100001",
       "01100101",
       "01100010",
       "01100000",
       "01100000",
       "01100010",
       "01100100",
       "01100011",
       "01100000",
       "01100000",
       "01010110",
       "01001100",
       "01001101",
       "01001000",
       "01000110",
       "01001100",
       "01001010",
       "00100111",
       "00010001",
       "00001110",
       "00001101",
       "00000111",
       "00001000",
       "00001111",
       "00100000",
       "01000111",
       "01011100",
       "01011010",
       "01011100",
       "01011100",
       "00111100",
       "00011001",
       "00001100",
       "00001001",
       "00001111",
       "00010101",
       "00001110",
       "00010011",
       "00010010",
       "00101011",
       "01001001",
       "01001100",
       "01001100",
       "01001011",
       "01011000",
       "01100001",
       "01100010",
       "01100100",
       "01100010",
       "01011111",
       "01100010",
       "01011101",
       "01100000",
       "01010110",
       "01010000",
       "01011001",
       "01011001",
       "01011100",
       "01100010",
       "01100101",
       "01100100",
       "01100001",
       "01100011",
       "01100100",
       "01100000",
       "01100000",
       "01100000",
       "01100001",
       "01011110",
       "01010100",
       "01001101",
       "01001011",
       "01001011",
       "01001111",
       "01010001",
       "01011010",
       "01011101",
       "01011101",
       "01011100",
       "01011101",
       "01010110",
       "01010010",
       "01001000",
       "01000001",
       "00111111",
       "00111101",
       "00100011",
       "00011100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00100100",
       "00010101",
       "00101001",
       "00011111",
       "00111111",
       "01000001",
       "01001010",
       "01011000",
       "01010111",
       "01001100",
       "01000011",
       "00111110",
       "00111000",
       "00011110",
       "00101000",
       "00110111",
       "00111011",
       "00111110",
       "00111110",
       "01000000",
       "01000101",
       "01001101",
       "01010010",
       "01011100",
       "01011111",
       "01011110",
       "01011110",
       "01011111",
       "01011110",
       "01100001",
       "01011110",
       "01100010",
       "01011000",
       "01010100",
       "01100100",
       "01100011",
       "01100011",
       "01100000",
       "01011110",
       "01011011",
       "01010001",
       "01001100",
       "01001100",
       "01000110",
       "01000011",
       "00111110",
       "01000011",
       "00111111",
       "00010111",
       "00010100",
       "00010001",
       "00010101",
       "00010001",
       "00010000",
       "00001101",
       "00001111",
       "00110011",
       "01000010",
       "01001001",
       "00101110",
       "00001011",
       "00010000",
       "00010010",
       "00011000",
       "00010100",
       "00010001",
       "00001010",
       "00001111",
       "00100100",
       "01001000",
       "01001000",
       "01001101",
       "01001110",
       "01010011",
       "01011000",
       "01011111",
       "01100110",
       "01100101",
       "01100011",
       "01100101",
       "01100010",
       "01100001",
       "01011110",
       "01011100",
       "01010110",
       "01011000",
       "01010110",
       "01010000",
       "01010001",
       "01011010",
       "01100000",
       "01100001",
       "01100000",
       "01100001",
       "01011110",
       "01100011",
       "01100000",
       "01100001",
       "01011100",
       "01100001",
       "01011101",
       "01011110",
       "01011101",
       "01011101",
       "01011111",
       "01011111",
       "01100000",
       "01100000",
       "01011100",
       "01011101",
       "01010011",
       "01010011",
       "01001000",
       "01000011",
       "00111101",
       "00111111",
       "00011110",
       "00011111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00100011",
       "00010010",
       "00101101",
       "00011110",
       "00111110",
       "01000000",
       "01001010",
       "01010100",
       "01010111",
       "01001000",
       "01000101",
       "00111101",
       "00111000",
       "00100000",
       "00010100",
       "00100011",
       "00110111",
       "00111010",
       "00111011",
       "01000100",
       "01001101",
       "01010011",
       "01011010",
       "01011110",
       "01011100",
       "01011000",
       "01010010",
       "01010000",
       "01010000",
       "01010010",
       "01010110",
       "01011011",
       "01010111",
       "01010111",
       "01100101",
       "01100000",
       "01100110",
       "01100011",
       "01100000",
       "01011011",
       "01011000",
       "01010011",
       "01001100",
       "01001111",
       "00111001",
       "00111010",
       "01000101",
       "01001010",
       "00101001",
       "00001110",
       "00010100",
       "00010010",
       "00010011",
       "00010001",
       "00011100",
       "00001101",
       "00101001",
       "00111100",
       "01000010",
       "00100010",
       "00010001",
       "00011000",
       "00010000",
       "00010000",
       "00001110",
       "00010010",
       "00010010",
       "00010100",
       "00111010",
       "01001110",
       "01001001",
       "01010000",
       "01010000",
       "01011010",
       "01011011",
       "01100010",
       "01100011",
       "01100011",
       "01100000",
       "01100111",
       "01100110",
       "01100100",
       "01010110",
       "01010011",
       "01011011",
       "01011010",
       "01011000",
       "01010100",
       "01010000",
       "01010100",
       "01011001",
       "01011111",
       "01011111",
       "01100001",
       "01100000",
       "01100001",
       "01011101",
       "01011101",
       "01010110",
       "01011110",
       "01011111",
       "01100010",
       "01100010",
       "01100011",
       "01100010",
       "01100100",
       "01100001",
       "01100000",
       "01011010",
       "01011011",
       "01010100",
       "01010100",
       "01000101",
       "01000011",
       "00111110",
       "01000000",
       "00010111",
       "00011111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010111",
       "00101101",
       "00011110",
       "00110000",
       "00110000",
       "01000100",
       "01000001",
       "01001011",
       "01010001",
       "01010101",
       "01000111",
       "01000001",
       "00111011",
       "00110110",
       "00011101",
       "00010001",
       "00101000",
       "00111101",
       "00111010",
       "00111111",
       "01001001",
       "01010101",
       "01010110",
       "01011000",
       "01011000",
       "01010001",
       "01001010",
       "00111110",
       "01000001",
       "01000000",
       "01000010",
       "01010010",
       "01010011",
       "01011011",
       "01100100",
       "01100011",
       "01100110",
       "01100110",
       "01100000",
       "01100011",
       "01100001",
       "01100001",
       "01010111",
       "01001111",
       "01010001",
       "00111111",
       "01000101",
       "01001000",
       "01001010",
       "00111001",
       "00010100",
       "00010111",
       "00010000",
       "00010100",
       "00010000",
       "00010011",
       "00001110",
       "00100101",
       "01000110",
       "01000101",
       "00100000",
       "00010010",
       "00010011",
       "00010010",
       "00010110",
       "00010011",
       "00011000",
       "00010100",
       "00100001",
       "01000111",
       "01001100",
       "01001101",
       "01001111",
       "01010110",
       "01011010",
       "01100011",
       "01100011",
       "01100011",
       "01100110",
       "01100110",
       "01100101",
       "01100101",
       "01100001",
       "01011100",
       "01001011",
       "01010000",
       "01011001",
       "01010001",
       "01010000",
       "01000110",
       "01000001",
       "01000101",
       "01000111",
       "01001110",
       "01011000",
       "01011010",
       "01011110",
       "01100000",
       "01011011",
       "01011001",
       "01011101",
       "01011101",
       "01100100",
       "01011101",
       "01011100",
       "01100000",
       "01100011",
       "01011100",
       "01100000",
       "01011001",
       "01011010",
       "01010111",
       "01010011",
       "01000111",
       "01000100",
       "00111010",
       "01000001",
       "00011110",
       "00100001",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00011100",
       "00101100",
       "00101100",
       "00110000",
       "00111110",
       "01000010",
       "01000100",
       "01001011",
       "01010111",
       "01010010",
       "01000101",
       "01000000",
       "00111011",
       "00101011",
       "00010110",
       "00011100",
       "00111100",
       "00111100",
       "00111111",
       "01000111",
       "01010011",
       "01010111",
       "01010100",
       "01010010",
       "01001011",
       "01000101",
       "01000010",
       "00111010",
       "00110011",
       "00110101",
       "00111100",
       "01001010",
       "01010101",
       "01010111",
       "01100101",
       "01100010",
       "01100111",
       "01100100",
       "01100011",
       "01100011",
       "01100011",
       "01100010",
       "01011101",
       "01010111",
       "01010000",
       "01001010",
       "01001100",
       "01001101",
       "01000111",
       "00111100",
       "00011111",
       "00010001",
       "00010000",
       "00010001",
       "00010101",
       "00010101",
       "00010001",
       "00011010",
       "00111110",
       "01001001",
       "00011111",
       "00010101",
       "00010101",
       "00010110",
       "00011000",
       "00010010",
       "00011000",
       "00010001",
       "00101111",
       "01001100",
       "01001101",
       "01010011",
       "01010011",
       "01010101",
       "01100101",
       "01100110",
       "01101001",
       "01100111",
       "01100111",
       "01100101",
       "01100111",
       "01100001",
       "01100000",
       "01100010",
       "01010111",
       "01001011",
       "01010011",
       "01000000",
       "00111111",
       "00111101",
       "00111100",
       "00110111",
       "00111000",
       "00111100",
       "01000001",
       "01000110",
       "01010000",
       "01010100",
       "01011101",
       "01011110",
       "01100010",
       "01011111",
       "01100101",
       "01100000",
       "01100000",
       "01011001",
       "01011110",
       "01011011",
       "01011110",
       "01011000",
       "01010101",
       "01010010",
       "01010001",
       "01000110",
       "01000100",
       "00110110",
       "00111110",
       "00011111",
       "00011001",
       "00010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00110110",
       "00101101",
       "00100101",
       "00101000",
       "00111010",
       "01000001",
       "00111111",
       "01001000",
       "01001111",
       "01010110",
       "01001101",
       "01000100",
       "00111110",
       "00110001",
       "00100001",
       "00010111",
       "00100110",
       "00111100",
       "00111100",
       "01001110",
       "01010010",
       "01010111",
       "01010100",
       "01010011",
       "01000101",
       "00111101",
       "00111011",
       "00111111",
       "00110001",
       "00101011",
       "00110111",
       "01000001",
       "01001010",
       "01011001",
       "01011011",
       "01100101",
       "01100011",
       "01100010",
       "01100001",
       "01100000",
       "01100001",
       "01101000",
       "01100010",
       "01100001",
       "01100100",
       "01011011",
       "01010000",
       "01001111",
       "01010011",
       "01001011",
       "01000011",
       "00101111",
       "00001110",
       "00010001",
       "00010010",
       "00010101",
       "00010001",
       "00010101",
       "00010110",
       "01000101",
       "01001011",
       "00100001",
       "00010001",
       "00010101",
       "00010001",
       "00010111",
       "00010001",
       "00011000",
       "00010110",
       "00111101",
       "01001010",
       "01010011",
       "01010011",
       "01010101",
       "01010111",
       "01101000",
       "01100101",
       "01101010",
       "01101010",
       "01101011",
       "01100111",
       "01101000",
       "01100100",
       "01100100",
       "01100000",
       "01011111",
       "01010010",
       "01001101",
       "00111101",
       "00111110",
       "00110000",
       "00111011",
       "00110111",
       "00111100",
       "00111010",
       "00110111",
       "00111001",
       "00111111",
       "01000000",
       "01001110",
       "01011010",
       "01100011",
       "01011100",
       "01100100",
       "01011111",
       "01100001",
       "01011000",
       "01011110",
       "01011100",
       "01011010",
       "01010001",
       "01010001",
       "01001110",
       "01001111",
       "01000101",
       "01000010",
       "00111000",
       "00111111",
       "00100100",
       "00010111",
       "00100100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00101101",
       "00101100",
       "00100111",
       "00100110",
       "00111100",
       "01000011",
       "01000001",
       "01001001",
       "01001111",
       "01010101",
       "01001100",
       "01000100",
       "00111011",
       "00110001",
       "00101011",
       "00100000",
       "00110000",
       "00111101",
       "00111110",
       "01010101",
       "01011001",
       "01011001",
       "01010010",
       "01001001",
       "00110111",
       "00111010",
       "00110111",
       "00101011",
       "00101000",
       "00111000",
       "00111110",
       "00111111",
       "01001101",
       "01011000",
       "01011111",
       "01101000",
       "01100000",
       "01100000",
       "01010111",
       "01011110",
       "01100001",
       "01100111",
       "01100111",
       "01100110",
       "01100110",
       "01100100",
       "01010110",
       "01010001",
       "01001101",
       "01001110",
       "01000110",
       "00111000",
       "00010100",
       "00010110",
       "00010001",
       "00010101",
       "00010101",
       "00011010",
       "00011001",
       "01000011",
       "01010011",
       "00100110",
       "00010000",
       "00010111",
       "00010110",
       "00011000",
       "00010110",
       "00010111",
       "00011110",
       "01001000",
       "01001111",
       "01010011",
       "01010100",
       "01011101",
       "01100110",
       "01100111",
       "01101000",
       "01101001",
       "01101001",
       "01101011",
       "01100110",
       "01101001",
       "01100100",
       "01100011",
       "01011110",
       "01011101",
       "01011010",
       "01001110",
       "01000000",
       "00111111",
       "00011110",
       "00011111",
       "00100111",
       "00110000",
       "00110100",
       "00110101",
       "00110011",
       "00111000",
       "00111010",
       "00111100",
       "01000101",
       "01010110",
       "01010111",
       "01100010",
       "01100000",
       "01011111",
       "01011111",
       "01011101",
       "01011001",
       "01010111",
       "01001001",
       "01001101",
       "01000111",
       "01001101",
       "01000101",
       "01000100",
       "00111101",
       "01000101",
       "00110000",
       "00011111",
       "00111100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00011011",
       "00100011",
       "00100000",
       "00101000",
       "00111101",
       "01001010",
       "01000001",
       "01001011",
       "01001111",
       "01010011",
       "01001001",
       "00111110",
       "00111110",
       "00111111",
       "00110101",
       "00101101",
       "00110011",
       "00111101",
       "00111101",
       "01010011",
       "01011001",
       "01011001",
       "01000111",
       "00111100",
       "00110110",
       "00110101",
       "00100010",
       "00100110",
       "00111000",
       "00111110",
       "01000001",
       "01000011",
       "01010000",
       "01010110",
       "01100000",
       "01100110",
       "01011010",
       "01011100",
       "01010011",
       "01011100",
       "01100000",
       "01100101",
       "01101010",
       "01101110",
       "01101010",
       "01101001",
       "01011110",
       "01011001",
       "01010001",
       "01010011",
       "01000110",
       "00111111",
       "00011110",
       "00010100",
       "00010001",
       "00010001",
       "00011000",
       "00010111",
       "00011101",
       "01000110",
       "01011001",
       "00110011",
       "00010111",
       "00011010",
       "00011000",
       "00011001",
       "00011001",
       "00010110",
       "00011100",
       "01001000",
       "01010011",
       "01010110",
       "01011010",
       "01101000",
       "01101011",
       "01101010",
       "01101000",
       "01101011",
       "01100110",
       "01101000",
       "01100011",
       "01100001",
       "01011100",
       "01011011",
       "01100100",
       "01011100",
       "01011010",
       "01001111",
       "01000100",
       "01000101",
       "00101110",
       "00011010",
       "00010101",
       "00010111",
       "00011111",
       "00100110",
       "00101010",
       "00101111",
       "00110010",
       "00111011",
       "00111011",
       "01000011",
       "01010000",
       "01011100",
       "01011111",
       "01100000",
       "01011111",
       "01100000",
       "01011001",
       "01010101",
       "01000101",
       "01000011",
       "01000001",
       "01001000",
       "01000100",
       "01000101",
       "00111101",
       "00111111",
       "00110110",
       "00101011",
       "00101011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00110100",
       "00101010",
       "00011011",
       "00011110",
       "00111010",
       "01000111",
       "01000010",
       "01001010",
       "01010001",
       "01010100",
       "01001100",
       "01000001",
       "00111111",
       "00111111",
       "00111001",
       "00111001",
       "00110101",
       "00111001",
       "01000000",
       "01010000",
       "01010110",
       "01001011",
       "00111110",
       "00111001",
       "00110001",
       "00011101",
       "00100010",
       "00110111",
       "00111111",
       "01000001",
       "01000001",
       "01000111",
       "01010100",
       "01011000",
       "01100011",
       "01100000",
       "01011010",
       "01011001",
       "01010100",
       "01010110",
       "01011011",
       "01100111",
       "01101000",
       "01101111",
       "01101010",
       "01100101",
       "01100001",
       "01100100",
       "01010110",
       "01010010",
       "01001000",
       "01000010",
       "00110100",
       "00010010",
       "00010101",
       "00010101",
       "00011011",
       "00011100",
       "00110001",
       "01011011",
       "01100000",
       "01000010",
       "00010101",
       "00011001",
       "00011000",
       "00010110",
       "00011001",
       "00010101",
       "00101000",
       "01001000",
       "01001001",
       "01011000",
       "01011011",
       "01100111",
       "01100110",
       "01101111",
       "01101100",
       "01101101",
       "01101000",
       "01100001",
       "01100001",
       "01011010",
       "01011001",
       "01010100",
       "01011110",
       "01011100",
       "01010001",
       "01010100",
       "01000011",
       "01001000",
       "00111000",
       "00011111",
       "00011000",
       "00010111",
       "00010011",
       "00010110",
       "00011110",
       "00100101",
       "00101010",
       "00110001",
       "00111000",
       "01000000",
       "01000101",
       "01001110",
       "01011010",
       "01011100",
       "01010111",
       "01100001",
       "01011001",
       "01001110",
       "01000111",
       "01000101",
       "01000001",
       "01000100",
       "01000000",
       "01000101",
       "00111100",
       "00111111",
       "00110101",
       "00101110",
       "00100111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00011100",
       "00001111",
       "00100100",
       "00101110",
       "01000101",
       "01000001",
       "01001011",
       "01001111",
       "01010110",
       "01001110",
       "01000111",
       "00111111",
       "00111100",
       "00111011",
       "00111011",
       "00111001",
       "00111011",
       "01000000",
       "01001110",
       "01010110",
       "01001000",
       "00111011",
       "00111100",
       "00011101",
       "00011001",
       "00111010",
       "00111101",
       "01000001",
       "01000010",
       "01001011",
       "01001101",
       "01010100",
       "01011111",
       "01100101",
       "01011101",
       "01011101",
       "01010111",
       "01010010",
       "01010100",
       "01010101",
       "01011100",
       "01100011",
       "01100110",
       "01100011",
       "01100101",
       "01101001",
       "01100111",
       "01100000",
       "01001100",
       "01001101",
       "00111111",
       "01000101",
       "00101000",
       "00010101",
       "00010101",
       "00010111",
       "00100101",
       "01001001",
       "01100101",
       "01100111",
       "01011011",
       "00101010",
       "00010011",
       "00010110",
       "00010101",
       "00010111",
       "00010111",
       "00110110",
       "01001100",
       "01001111",
       "01011101",
       "01100010",
       "01101000",
       "01100111",
       "01101100",
       "01101011",
       "01101111",
       "01100110",
       "01011011",
       "01011010",
       "01010111",
       "01010111",
       "01010110",
       "01011000",
       "01011111",
       "01010011",
       "01010011",
       "01000110",
       "01000110",
       "00110111",
       "00100000",
       "00011010",
       "00010111",
       "00011001",
       "00001111",
       "00010110",
       "00011110",
       "00100000",
       "00100101",
       "00100110",
       "00110100",
       "00111111",
       "01001000",
       "01001111",
       "01010111",
       "01011010",
       "01010110",
       "01011001",
       "01010001",
       "01001001",
       "01001000",
       "01000001",
       "01000100",
       "00111110",
       "01000101",
       "00111010",
       "01000100",
       "00111000",
       "00101110",
       "00001110",
       "00010100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010011",
       "00010010",
       "00110110",
       "00101100",
       "01001010",
       "01000001",
       "01000111",
       "01001101",
       "01010101",
       "01001011",
       "01001110",
       "01000111",
       "01000011",
       "01000001",
       "00111101",
       "00111101",
       "00111111",
       "01000011",
       "01010010",
       "01010011",
       "01000100",
       "00111110",
       "00110010",
       "00010100",
       "00110110",
       "00111101",
       "00111110",
       "00111111",
       "01000011",
       "01001110",
       "01010001",
       "01010111",
       "01100000",
       "01011100",
       "01011011",
       "01011010",
       "01010101",
       "01010001",
       "01010100",
       "01010011",
       "01010100",
       "01010001",
       "01100000",
       "01101010",
       "01101001",
       "01101011",
       "01101000",
       "01100111",
       "01011000",
       "01010011",
       "01001011",
       "00111110",
       "00111111",
       "00011111",
       "00010110",
       "00100000",
       "00110000",
       "01001111",
       "01101010",
       "01100011",
       "01100100",
       "01000111",
       "00100010",
       "00100001",
       "00011010",
       "00011010",
       "00011001",
       "00111100",
       "01010110",
       "01011001",
       "01100101",
       "01100010",
       "01101011",
       "01100111",
       "01101100",
       "01101010",
       "01101000",
       "01011111",
       "01011010",
       "01010101",
       "01010010",
       "01010101",
       "01011001",
       "01010110",
       "01011101",
       "01011001",
       "01010001",
       "01001011",
       "01000100",
       "00111110",
       "00101101",
       "00011001",
       "00011010",
       "00011101",
       "00010111",
       "00001110",
       "00011110",
       "00011010",
       "00011110",
       "00011011",
       "00100111",
       "00110111",
       "01000010",
       "01000101",
       "01001111",
       "01011001",
       "01011001",
       "01010101",
       "01011010",
       "01001100",
       "01000101",
       "01000000",
       "01000001",
       "00111100",
       "01000010",
       "00111111",
       "01000011",
       "00111101",
       "00101110",
       "00010011",
       "00011010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001110",
       "00111001",
       "00100101",
       "01000111",
       "01000011",
       "01000101",
       "01001011",
       "01001111",
       "01010000",
       "01010010",
       "01010011",
       "01001001",
       "01000100",
       "00111111",
       "01000000",
       "01000100",
       "01001010",
       "01011000",
       "01010100",
       "00111110",
       "01000000",
       "00100110",
       "00100111",
       "01000000",
       "00110111",
       "00111110",
       "01000011",
       "01001101",
       "01010001",
       "01011100",
       "01010111",
       "01011111",
       "01011001",
       "01010111",
       "01010111",
       "01010100",
       "01010110",
       "01010100",
       "01010111",
       "01010001",
       "01000011",
       "01011101",
       "01100110",
       "01101001",
       "01101001",
       "01101011",
       "01101001",
       "01101001",
       "01011001",
       "01010001",
       "00111010",
       "00111010",
       "00101000",
       "00011000",
       "00100001",
       "00101100",
       "01010111",
       "01101101",
       "01101000",
       "01011111",
       "01000010",
       "00110010",
       "00101000",
       "00011100",
       "00100000",
       "00011010",
       "01000100",
       "01011111",
       "01100000",
       "01101001",
       "01100110",
       "01101101",
       "01101001",
       "01110010",
       "01101101",
       "01101001",
       "01011010",
       "01010101",
       "01010011",
       "01010000",
       "01010001",
       "01011000",
       "01010100",
       "01011000",
       "01011001",
       "01010001",
       "01001000",
       "01000100",
       "01000000",
       "00110010",
       "00101010",
       "00110100",
       "00110010",
       "00101111",
       "00010100",
       "00010010",
       "00011001",
       "00010100",
       "00011001",
       "00100110",
       "00110111",
       "00111110",
       "01000010",
       "01000110",
       "01001110",
       "01011010",
       "01010110",
       "01010111",
       "01010110",
       "01001011",
       "01000010",
       "01000100",
       "00111010",
       "01000000",
       "00111111",
       "01000010",
       "00111101",
       "00101110",
       "00011010",
       "00011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001010",
       "00001101",
       "00111011",
       "00100100",
       "00111000",
       "01000001",
       "01000011",
       "00111111",
       "01000101",
       "01000100",
       "01001101",
       "01001110",
       "01001101",
       "01001000",
       "01000100",
       "01000010",
       "01001001",
       "01010001",
       "01011000",
       "01010011",
       "01000000",
       "00111101",
       "00100010",
       "00101101",
       "00111101",
       "00111011",
       "01000010",
       "01001011",
       "01010011",
       "01010111",
       "01010111",
       "01010011",
       "01100011",
       "01011001",
       "01010101",
       "01010101",
       "01010011",
       "01010100",
       "01010101",
       "01010101",
       "01001011",
       "01001101",
       "01011011",
       "01100100",
       "01101001",
       "01101010",
       "01101100",
       "01101011",
       "01101011",
       "01100111",
       "01010110",
       "01001001",
       "00111111",
       "00110000",
       "00100110",
       "00011001",
       "00100000",
       "01000111",
       "01101100",
       "01101101",
       "01101111",
       "01001111",
       "00110111",
       "00100100",
       "00100011",
       "00011100",
       "00100101",
       "01010101",
       "01101000",
       "01101001",
       "01101010",
       "01101010",
       "01101101",
       "01101001",
       "01101101",
       "01101001",
       "01101000",
       "01011100",
       "01010001",
       "01010011",
       "01010110",
       "01010010",
       "01010110",
       "01010111",
       "01010111",
       "01011010",
       "01010100",
       "01001010",
       "01001000",
       "01000001",
       "00111011",
       "00111001",
       "01000011",
       "01000001",
       "01000011",
       "00110010",
       "00001111",
       "00001111",
       "00001101",
       "00011000",
       "00101001",
       "00111101",
       "01000011",
       "01000011",
       "01000100",
       "01000101",
       "01010001",
       "01010110",
       "01010111",
       "01011000",
       "01010101",
       "01000111",
       "01000101",
       "00111101",
       "01000101",
       "00111001",
       "00111110",
       "00101111",
       "00101011",
       "00010110",
       "00010100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010011",
       "00111110",
       "00100110",
       "00011010",
       "00110011",
       "01000011",
       "01000000",
       "00111110",
       "00111010",
       "01000001",
       "00111100",
       "01000011",
       "01000110",
       "01001011",
       "01000000",
       "01000111",
       "01010011",
       "01011000",
       "01000111",
       "01000001",
       "00111011",
       "00011011",
       "00110010",
       "01000010",
       "00111011",
       "00111110",
       "01001000",
       "01010010",
       "01010100",
       "01010010",
       "01010100",
       "01011111",
       "01010110",
       "01011000",
       "01010101",
       "01010011",
       "01010110",
       "01011010",
       "01010000",
       "01010101",
       "01011011",
       "01100011",
       "01100111",
       "01100110",
       "01101001",
       "01101101",
       "01101110",
       "01101100",
       "01101011",
       "01101001",
       "01011110",
       "01001111",
       "01000000",
       "00110011",
       "00100101",
       "00100001",
       "00101110",
       "01010110",
       "01011000",
       "01100100",
       "01001000",
       "00110100",
       "00011111",
       "00101000",
       "00101101",
       "01000011",
       "01100001",
       "01101011",
       "01101000",
       "01101010",
       "01101100",
       "01101101",
       "01101010",
       "01101000",
       "01101001",
       "01100011",
       "01011100",
       "01010011",
       "01001100",
       "01011000",
       "01010111",
       "01010001",
       "01010110",
       "01010011",
       "01011001",
       "01010111",
       "01010000",
       "01001101",
       "01000001",
       "01000011",
       "01000100",
       "01000100",
       "00111110",
       "01000010",
       "01000100",
       "00101001",
       "00001111",
       "00001111",
       "00010101",
       "00110010",
       "00111010",
       "01000110",
       "01000011",
       "01000111",
       "01000110",
       "01001110",
       "01001111",
       "01011011",
       "01010100",
       "01011000",
       "01001111",
       "01000111",
       "00111111",
       "01000011",
       "00110011",
       "00111010",
       "00011111",
       "00100010",
       "00010110",
       "00010111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00100010",
       "00111100",
       "00110101",
       "00100100",
       "00011100",
       "00110010",
       "00101100",
       "00111011",
       "00110110",
       "01000001",
       "00111011",
       "00111111",
       "00111011",
       "01000011",
       "00111111",
       "01000111",
       "01010011",
       "01010011",
       "01000000",
       "00111101",
       "00110111",
       "00011001",
       "00110111",
       "01000001",
       "00111101",
       "00111111",
       "01000010",
       "01001100",
       "01010010",
       "01001010",
       "01010001",
       "01011111",
       "01010101",
       "01011000",
       "01011000",
       "01011001",
       "01010010",
       "01010000",
       "01010011",
       "01011100",
       "01100000",
       "01100101",
       "01011110",
       "01100001",
       "01100111",
       "01101101",
       "01110011",
       "01101011",
       "01101001",
       "01101010",
       "01100001",
       "01011100",
       "01001111",
       "00111110",
       "00011010",
       "00100000",
       "00100010",
       "00111000",
       "00111111",
       "00111001",
       "01000001",
       "00100111",
       "00011010",
       "00101000",
       "01001011",
       "01011111",
       "01100110",
       "01101001",
       "01101010",
       "01101011",
       "01101101",
       "01101010",
       "01101000",
       "01101001",
       "01100111",
       "01100011",
       "01011110",
       "01011011",
       "01010011",
       "01010001",
       "01010110",
       "01001111",
       "01010110",
       "01010100",
       "01010100",
       "01010111",
       "01010100",
       "01010100",
       "01001100",
       "01000111",
       "01001011",
       "01001001",
       "01000011",
       "00111100",
       "00111111",
       "00111100",
       "00011000",
       "00010001",
       "00010110",
       "00110001",
       "00111110",
       "01000100",
       "01000100",
       "01000010",
       "01000100",
       "01001010",
       "01001110",
       "01010101",
       "01010101",
       "01010010",
       "01001110",
       "01001000",
       "00111101",
       "01000001",
       "00110000",
       "00101111",
       "00010110",
       "00100011",
       "00011110",
       "00010100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00101001",
       "00110101",
       "00111000",
       "00100101",
       "00001111",
       "00100000",
       "00011001",
       "00101100",
       "00101101",
       "00110010",
       "00111000",
       "01000011",
       "00111101",
       "00111011",
       "00111101",
       "01001001",
       "01001101",
       "01001011",
       "00111110",
       "00111111",
       "00110000",
       "00100001",
       "00111000",
       "00111111",
       "01000000",
       "00111110",
       "00111110",
       "01001111",
       "01001011",
       "01000011",
       "01010011",
       "01011101",
       "01010001",
       "01010100",
       "01011000",
       "01010110",
       "01000101",
       "01010011",
       "01011001",
       "01011111",
       "01100001",
       "01100010",
       "01011110",
       "01011111",
       "01100000",
       "01100101",
       "01101100",
       "01101101",
       "01101011",
       "01101010",
       "01100010",
       "01100011",
       "01011101",
       "01010101",
       "00100111",
       "00011111",
       "00011001",
       "00011100",
       "00100000",
       "00011000",
       "00110101",
       "00011101",
       "00100101",
       "00111110",
       "01011010",
       "01101101",
       "01101000",
       "01101001",
       "01100110",
       "01101011",
       "01101011",
       "01101001",
       "01100010",
       "01100011",
       "01100000",
       "01100000",
       "01100010",
       "01011100",
       "01011100",
       "01010111",
       "01011010",
       "01011001",
       "01010111",
       "01010101",
       "01010100",
       "01011001",
       "01010100",
       "01010001",
       "01010010",
       "01010110",
       "01010001",
       "01010010",
       "01000111",
       "01000010",
       "00111110",
       "00111010",
       "00100101",
       "00010000",
       "00010110",
       "00101011",
       "00111101",
       "00111100",
       "01000001",
       "00111110",
       "01000010",
       "01001001",
       "01010010",
       "01010110",
       "01011001",
       "01010011",
       "01010000",
       "01001010",
       "00111100",
       "00111110",
       "00110010",
       "00011110",
       "00001110",
       "00101100",
       "00100100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001000",
       "00101101",
       "00011011",
       "00011110",
       "00011001",
       "00101011",
       "00110000",
       "00101100",
       "00101101",
       "00101000",
       "00011110",
       "00011011",
       "00101100",
       "00110110",
       "00111110",
       "00111010",
       "01000000",
       "01000110",
       "01000111",
       "00111011",
       "00110110",
       "00100100",
       "00101001",
       "00110111",
       "00111101",
       "01000000",
       "01000000",
       "01000001",
       "01010010",
       "00111100",
       "01001001",
       "01011111",
       "01011000",
       "01010101",
       "01010100",
       "01011001",
       "01010100",
       "01001010",
       "01011110",
       "01011101",
       "01100001",
       "01100100",
       "01100001",
       "01011111",
       "01100000",
       "01100001",
       "01100001",
       "01101000",
       "01110000",
       "01101010",
       "01101010",
       "01100010",
       "01100110",
       "01100101",
       "01100011",
       "01001111",
       "00101000",
       "00100001",
       "00011001",
       "00010011",
       "00010100",
       "00100001",
       "00100000",
       "00111101",
       "01100100",
       "01011111",
       "01101011",
       "01100111",
       "01100111",
       "01101000",
       "01101100",
       "01101100",
       "01100110",
       "01011111",
       "01011100",
       "01100000",
       "01011111",
       "01100000",
       "01100001",
       "01011110",
       "01011100",
       "01011011",
       "01011010",
       "01010110",
       "01010001",
       "01010101",
       "01010111",
       "01010011",
       "01001111",
       "01010001",
       "01010100",
       "01001011",
       "01001011",
       "01000110",
       "01000101",
       "00111111",
       "00111010",
       "00101110",
       "00010000",
       "00011010",
       "00011011",
       "00110001",
       "01000000",
       "00111101",
       "00110110",
       "00111101",
       "01000010",
       "01001101",
       "01010000",
       "01010010",
       "01001111",
       "01001101",
       "01001001",
       "01000001",
       "00111100",
       "00110111",
       "00001101",
       "00010011",
       "00101000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000110",
       "00100110",
       "00001111",
       "00100110",
       "00111001",
       "01000100",
       "00111110",
       "00111101",
       "00111101",
       "00110110",
       "00101100",
       "00011001",
       "00011100",
       "00100011",
       "00101110",
       "00111100",
       "00111100",
       "01000000",
       "00111011",
       "01000000",
       "00100011",
       "00011101",
       "00100011",
       "00110001",
       "00111111",
       "00111110",
       "01000001",
       "01000110",
       "00111110",
       "00100100",
       "01000111",
       "01011001",
       "01011001",
       "01011000",
       "01010111",
       "01011010",
       "01010110",
       "01010010",
       "01011001",
       "01100000",
       "01100011",
       "01100010",
       "01100010",
       "01100011",
       "01100001",
       "01100101",
       "01100100",
       "01101011",
       "01101111",
       "01101101",
       "01101110",
       "01100101",
       "01101001",
       "01100111",
       "01011111",
       "01100001",
       "00110011",
       "00011101",
       "00100010",
       "00010100",
       "00011011",
       "00100011",
       "00101101",
       "01010011",
       "01100111",
       "01100011",
       "01101001",
       "01101100",
       "01101001",
       "01101100",
       "01101101",
       "01101110",
       "01100101",
       "01100000",
       "01011101",
       "01100000",
       "01011110",
       "01011101",
       "01100100",
       "01100001",
       "01011101",
       "01010111",
       "01010101",
       "01011001",
       "01010010",
       "01010010",
       "01010110",
       "01011000",
       "01001010",
       "01001011",
       "01001010",
       "01000011",
       "00111111",
       "00111100",
       "00111111",
       "00111110",
       "00111101",
       "00110100",
       "00010010",
       "00011001",
       "00010111",
       "00011001",
       "00110010",
       "01000000",
       "00111010",
       "00111111",
       "00111100",
       "01000100",
       "01000101",
       "01000101",
       "00111110",
       "01000000",
       "00111110",
       "01000001",
       "01000000",
       "00101110",
       "00000101",
       "00011100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001100",
       "00011100",
       "00100001",
       "01000010",
       "01000100",
       "01000110",
       "01000001",
       "01000101",
       "01000001",
       "01000001",
       "01000001",
       "00110010",
       "00100001",
       "00011100",
       "00010110",
       "00101010",
       "00111101",
       "01000100",
       "01000000",
       "01000100",
       "00011101",
       "00010111",
       "00011110",
       "00110011",
       "00111101",
       "01000000",
       "01000100",
       "01001110",
       "00111010",
       "00101100",
       "01001011",
       "01010101",
       "01010111",
       "01010000",
       "01010100",
       "01011000",
       "01010010",
       "01010100",
       "01011010",
       "01011111",
       "01100011",
       "01100101",
       "01100110",
       "01100111",
       "01101001",
       "01100101",
       "01100100",
       "01101000",
       "01101110",
       "01101011",
       "01101011",
       "01101000",
       "01101000",
       "01100110",
       "01011111",
       "01011110",
       "00111101",
       "00011010",
       "00011101",
       "00010010",
       "00011001",
       "00011101",
       "00111000",
       "01100001",
       "01100010",
       "01100110",
       "01101001",
       "01101011",
       "01101101",
       "01101100",
       "01101101",
       "01101011",
       "01101001",
       "01100111",
       "01100010",
       "01100110",
       "01100010",
       "01100001",
       "01011110",
       "01100101",
       "01100011",
       "01011010",
       "01011001",
       "01011001",
       "01001111",
       "01010001",
       "01010011",
       "01011001",
       "01001000",
       "01000110",
       "01000111",
       "01000100",
       "00111111",
       "00111010",
       "00111011",
       "00111001",
       "00111000",
       "00101000",
       "00010010",
       "00010100",
       "00011101",
       "00001111",
       "00010110",
       "00101001",
       "00110000",
       "00111011",
       "00111010",
       "00111110",
       "00111101",
       "00111111",
       "00111101",
       "01000001",
       "00111001",
       "00111010",
       "00110110",
       "00010001",
       "00000100",
       "00101001",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010000",
       "00010110",
       "00100011",
       "00110101",
       "01000110",
       "01000011",
       "01001010",
       "01000111",
       "01001100",
       "01000111",
       "01000000",
       "01000100",
       "00111110",
       "00111000",
       "00110000",
       "00101011",
       "00100011",
       "00101100",
       "00110110",
       "00111000",
       "00100111",
       "00011101",
       "00010011",
       "00011010",
       "00111000",
       "00111110",
       "01000011",
       "01000111",
       "01001111",
       "01001011",
       "00111110",
       "01001110",
       "01011000",
       "01010110",
       "01001111",
       "01010101",
       "01010100",
       "01010111",
       "01011000",
       "01011110",
       "01011101",
       "01100000",
       "01100101",
       "01101001",
       "01101001",
       "01101001",
       "01100000",
       "01100000",
       "01100101",
       "01101000",
       "01101011",
       "01101100",
       "01101010",
       "01100111",
       "01100100",
       "01011101",
       "01010110",
       "01000101",
       "00011100",
       "00011010",
       "00010010",
       "00011001",
       "00011011",
       "00110101",
       "01011100",
       "01100000",
       "01100011",
       "01100110",
       "01101100",
       "01110001",
       "01101011",
       "01101110",
       "01101001",
       "01100100",
       "01100110",
       "01100011",
       "01100011",
       "01100011",
       "01100110",
       "01100001",
       "01100011",
       "01100000",
       "01011100",
       "01011000",
       "01010100",
       "01001101",
       "01010001",
       "01010010",
       "01010110",
       "01001101",
       "01010000",
       "01000101",
       "01000001",
       "01000001",
       "00111100",
       "00111001",
       "00110000",
       "00100011",
       "00010111",
       "00010000",
       "00010011",
       "00010111",
       "00010111",
       "00010011",
       "00010111",
       "00011000",
       "00100111",
       "00100101",
       "00100101",
       "00100101",
       "00101010",
       "00101101",
       "00110011",
       "00101101",
       "00100111",
       "00011011",
       "00010010",
       "00001110",
       "00011111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001100",
       "00010101",
       "00110100",
       "00111100",
       "00111110",
       "01000100",
       "01001010",
       "01001111",
       "01010110",
       "01010011",
       "01001100",
       "01000111",
       "01000011",
       "00111111",
       "01000000",
       "00111111",
       "00111100",
       "00100110",
       "00011010",
       "00011111",
       "00010010",
       "00010110",
       "00010011",
       "00010101",
       "00111001",
       "00111111",
       "01000001",
       "01000010",
       "01000111",
       "01010001",
       "01000110",
       "01010010",
       "01010010",
       "01011011",
       "01010000",
       "01010101",
       "01001000",
       "01010101",
       "01011101",
       "01100000",
       "01100000",
       "01100001",
       "01100000",
       "01101001",
       "01100110",
       "01100010",
       "01100011",
       "01100011",
       "01100100",
       "01100111",
       "01101100",
       "01110000",
       "01101110",
       "01101000",
       "01100101",
       "01011100",
       "01010001",
       "01001000",
       "00100001",
       "00011001",
       "00010100",
       "00010110",
       "00011000",
       "00110000",
       "01010010",
       "01010111",
       "01100001",
       "01100110",
       "01101111",
       "01101101",
       "01101111",
       "01101110",
       "01101000",
       "01100101",
       "01100001",
       "01100100",
       "01100001",
       "01100111",
       "01100110",
       "01100100",
       "01100010",
       "01100101",
       "01011011",
       "01010111",
       "01010010",
       "01010001",
       "01010011",
       "01010010",
       "01010100",
       "01001101",
       "01001111",
       "01001011",
       "01000110",
       "01000100",
       "00111110",
       "01000000",
       "00101011",
       "00011000",
       "00010100",
       "00001011",
       "00010001",
       "00010001",
       "00011100",
       "00100001",
       "00011111",
       "00011010",
       "00011100",
       "00011000",
       "00011011",
       "00011001",
       "00011001",
       "00010110",
       "00011101",
       "00011101",
       "00011110",
       "00011000",
       "00010110",
       "00010000",
       "00010011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010100",
       "00011011",
       "01000000",
       "00111100",
       "00111100",
       "01000011",
       "01001100",
       "01010110",
       "01011010",
       "01011001",
       "01010110",
       "01011000",
       "01010001",
       "01000101",
       "00111111",
       "00111110",
       "01000010",
       "00111100",
       "00101101",
       "00011110",
       "00010010",
       "00010011",
       "00001100",
       "00010101",
       "00100010",
       "00110101",
       "01000001",
       "01000010",
       "01000110",
       "01010010",
       "01001110",
       "01010001",
       "01001101",
       "01011000",
       "01010010",
       "01010001",
       "01000000",
       "01001100",
       "01011100",
       "01100010",
       "01100010",
       "01100001",
       "01100111",
       "01101010",
       "01100101",
       "01100001",
       "01100010",
       "01100011",
       "01100011",
       "01101000",
       "01100111",
       "01110000",
       "01110000",
       "01100111",
       "01100101",
       "01011110",
       "01010101",
       "01010010",
       "00101001",
       "00011000",
       "00011000",
       "00011001",
       "00010111",
       "00110001",
       "01010110",
       "01010100",
       "01011111",
       "01100101",
       "01101100",
       "01101101",
       "01110000",
       "01101011",
       "01100111",
       "01100110",
       "01011111",
       "01100100",
       "01100100",
       "01100101",
       "01100101",
       "01100011",
       "01100001",
       "01100011",
       "01011001",
       "01010111",
       "01010111",
       "01010101",
       "01010000",
       "01010100",
       "01010010",
       "01001101",
       "01010011",
       "01010011",
       "01001000",
       "01000110",
       "00111101",
       "00111110",
       "00101100",
       "00011101",
       "00011011",
       "00001110",
       "00010010",
       "00011011",
       "00100010",
       "00011111",
       "00011111",
       "00011011",
       "00011010",
       "00011010",
       "00100001",
       "00011110",
       "00100011",
       "00100000",
       "00100100",
       "00100110",
       "00101011",
       "00101010",
       "00100011",
       "00010100",
       "00010000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010101",
       "00011110",
       "00111101",
       "00111000",
       "00111011",
       "01000001",
       "01001001",
       "01010001",
       "01010010",
       "01010000",
       "01001111",
       "01010000",
       "01001100",
       "01010111",
       "01001010",
       "01000100",
       "00111110",
       "01000001",
       "01000000",
       "00101111",
       "00001111",
       "00010101",
       "00001010",
       "00010110",
       "00011101",
       "00111000",
       "01000001",
       "01000011",
       "01001000",
       "01010101",
       "01010011",
       "01010010",
       "01001010",
       "01010100",
       "01011001",
       "01001111",
       "01001001",
       "01010110",
       "01011000",
       "01100001",
       "01011110",
       "01011111",
       "01100011",
       "01100111",
       "01100101",
       "01100010",
       "01100001",
       "01100101",
       "01100011",
       "01101011",
       "01100101",
       "01101110",
       "01110000",
       "01100101",
       "01100010",
       "01011100",
       "01010010",
       "01011000",
       "00110011",
       "00011011",
       "00011100",
       "00011001",
       "00010110",
       "00110001",
       "01011000",
       "01010100",
       "01100001",
       "01100110",
       "01101100",
       "01110001",
       "01110011",
       "01101100",
       "01101010",
       "01100101",
       "01100000",
       "01011111",
       "01100101",
       "01100001",
       "01100011",
       "01100001",
       "01011110",
       "01011110",
       "01011100",
       "01011010",
       "01011001",
       "01010110",
       "01010010",
       "01001100",
       "01001001",
       "01001100",
       "01010010",
       "01010011",
       "01001010",
       "01000100",
       "00111110",
       "01000000",
       "00101011",
       "00010101",
       "00010100",
       "00010110",
       "00010000",
       "00010101",
       "00010111",
       "00011111",
       "00101000",
       "00100101",
       "00100011",
       "00011101",
       "00011011",
       "00011110",
       "00100100",
       "00101110",
       "00110101",
       "00111001",
       "00110110",
       "00111011",
       "00110101",
       "00110001",
       "00010110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010000",
       "00000110",
       "00100110",
       "00110001",
       "00111111",
       "00111001",
       "01000010",
       "00111111",
       "01001010",
       "01000011",
       "01000101",
       "01000010",
       "01000000",
       "00111101",
       "01011010",
       "01011000",
       "01001111",
       "01001000",
       "01000011",
       "00111110",
       "00111011",
       "00010101",
       "00010010",
       "00010001",
       "00011010",
       "00101101",
       "01000100",
       "01000001",
       "01001001",
       "01001110",
       "01010111",
       "01011011",
       "01010101",
       "01001100",
       "01001110",
       "01000111",
       "01010100",
       "01010001",
       "01011010",
       "01010101",
       "01011010",
       "01100010",
       "01100110",
       "01100011",
       "01101100",
       "01101000",
       "01100101",
       "01100101",
       "01101011",
       "01100100",
       "01101100",
       "01100110",
       "01101010",
       "01101100",
       "01100100",
       "01011111",
       "01100010",
       "01010010",
       "01011010",
       "01000101",
       "00100011",
       "00010110",
       "00010110",
       "00011000",
       "00110110",
       "01010011",
       "01011000",
       "01100010",
       "01101000",
       "01101111",
       "01110000",
       "01110100",
       "01110000",
       "01101100",
       "01101100",
       "01101001",
       "01100100",
       "01100110",
       "01100010",
       "01100011",
       "01100010",
       "01100000",
       "01011110",
       "01011110",
       "01011000",
       "01011000",
       "01010000",
       "01010011",
       "01001110",
       "01000101",
       "01001110",
       "01001110",
       "01001100",
       "01001000",
       "01000111",
       "00111110",
       "00111111",
       "00101111",
       "00010110",
       "00010000",
       "00010001",
       "00001110",
       "00010011",
       "00101001",
       "00111010",
       "00111101",
       "00111001",
       "00110010",
       "00101011",
       "00100000",
       "00011110",
       "00100111",
       "00111001",
       "00111111",
       "01000000",
       "00111001",
       "00111001",
       "00110111",
       "00111111",
       "00101100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00100001",
       "00010000",
       "00110111",
       "00100100",
       "01000000",
       "00111010",
       "01000000",
       "00111011",
       "00111111",
       "00111010",
       "00111100",
       "00111010",
       "00111110",
       "00111111",
       "01001011",
       "01010111",
       "01010111",
       "01010100",
       "01000111",
       "01000100",
       "00111011",
       "00010110",
       "00010010",
       "00010101",
       "00010110",
       "00100011",
       "01000010",
       "01000100",
       "01001000",
       "01001011",
       "01011000",
       "01011111",
       "01011000",
       "01001101",
       "01000000",
       "00110001",
       "01010110",
       "01010011",
       "01010111",
       "01010001",
       "01011001",
       "01010010",
       "01001111",
       "01001010",
       "01100101",
       "01100111",
       "01100111",
       "01100001",
       "01100011",
       "01100100",
       "01101011",
       "01100111",
       "01101011",
       "01101101",
       "01101000",
       "01100100",
       "01011111",
       "01011100",
       "01011000",
       "01001001",
       "00101010",
       "00010101",
       "00011001",
       "00011010",
       "00111111",
       "01010011",
       "01010111",
       "01011110",
       "01101000",
       "01101111",
       "01101100",
       "01101101",
       "01101100",
       "01110000",
       "01110000",
       "01101110",
       "01100110",
       "01100110",
       "01100100",
       "01100101",
       "01100100",
       "01100100",
       "01011101",
       "01100010",
       "01011101",
       "01011000",
       "01001110",
       "01001110",
       "01010001",
       "01001001",
       "01001110",
       "01001100",
       "01010000",
       "01000100",
       "01000001",
       "00111000",
       "00101011",
       "00101001",
       "00010111",
       "00011000",
       "00010101",
       "00001110",
       "00100011",
       "01000100",
       "01000011",
       "01000001",
       "00111110",
       "01000000",
       "01000000",
       "00110110",
       "00101100",
       "00111011",
       "00111101",
       "00111101",
       "00111001",
       "00111011",
       "00111000",
       "00111011",
       "00111001",
       "00110111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00110001",
       "00001101",
       "00110100",
       "00100110",
       "00111110",
       "00111010",
       "00111111",
       "00111010",
       "00111101",
       "00111100",
       "00111111",
       "00111010",
       "00111001",
       "00110101",
       "00111010",
       "01001101",
       "01011011",
       "01011001",
       "01001100",
       "01000100",
       "00111000",
       "00010101",
       "00010101",
       "00001101",
       "00010111",
       "00010111",
       "00111011",
       "01000001",
       "01000100",
       "01001000",
       "01011110",
       "01100001",
       "01011101",
       "01010011",
       "01001111",
       "00111100",
       "01001010",
       "01010010",
       "01011001",
       "01011010",
       "01100000",
       "01001000",
       "00101001",
       "00101110",
       "01010010",
       "01011101",
       "01100001",
       "01101000",
       "01100101",
       "01100111",
       "01100101",
       "01101001",
       "01100111",
       "01101000",
       "01101100",
       "01100111",
       "01011010",
       "01011101",
       "01011000",
       "01010011",
       "00110010",
       "00011000",
       "00011010",
       "00011100",
       "01000110",
       "01010100",
       "01010101",
       "01011011",
       "01100111",
       "01110000",
       "01101101",
       "01101101",
       "01101010",
       "01101100",
       "01101101",
       "01110000",
       "01100111",
       "01100110",
       "01100111",
       "01100101",
       "01100110",
       "01100100",
       "01100100",
       "01100000",
       "01010110",
       "01011010",
       "01001011",
       "01001101",
       "01010100",
       "01001100",
       "01001010",
       "01010001",
       "01010010",
       "01000101",
       "01000001",
       "00111110",
       "00100110",
       "00011110",
       "00100001",
       "00110001",
       "00011111",
       "00001100",
       "00110000",
       "01000100",
       "00111101",
       "01000100",
       "01000011",
       "01000101",
       "01000100",
       "00111111",
       "00111100",
       "00111110",
       "00111100",
       "01000001",
       "01000110",
       "01001001",
       "01000111",
       "01000011",
       "00110010",
       "00110101",
       "00010001",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010011",
       "00110000",
       "00010111",
       "01001000",
       "00111001",
       "01000011",
       "00111110",
       "01000110",
       "01000010",
       "01000101",
       "00111001",
       "00011111",
       "00101100",
       "01000011",
       "01000011",
       "01010111",
       "01010111",
       "01010001",
       "01000010",
       "00110001",
       "00010011",
       "00011001",
       "00001111",
       "00010110",
       "00010100",
       "00111000",
       "00111111",
       "01000100",
       "01010001",
       "01100000",
       "01011010",
       "01100001",
       "01011101",
       "01100011",
       "01010111",
       "01010011",
       "01000101",
       "01001111",
       "01101000",
       "01100101",
       "01010100",
       "01000001",
       "01001001",
       "01010011",
       "01010110",
       "01011000",
       "01011101",
       "01100011",
       "01101001",
       "01100011",
       "01100110",
       "01101001",
       "01100101",
       "01100111",
       "01101000",
       "01011100",
       "01011101",
       "01011010",
       "01011011",
       "00111000",
       "00011010",
       "00011110",
       "00100000",
       "01001001",
       "01010101",
       "01011011",
       "01100001",
       "01100110",
       "01101010",
       "01101000",
       "01101010",
       "01101101",
       "01101110",
       "01110000",
       "01110011",
       "01110000",
       "01101100",
       "01100011",
       "01011100",
       "01100010",
       "01011010",
       "01010110",
       "01001011",
       "01000011",
       "01001001",
       "01001000",
       "01001111",
       "01011011",
       "01010011",
       "01001100",
       "01010100",
       "01010010",
       "01001100",
       "01000101",
       "01000011",
       "00111001",
       "00110100",
       "00110110",
       "00110000",
       "00010000",
       "00010001",
       "00101101",
       "01000101",
       "01000000",
       "01001011",
       "01001101",
       "01010001",
       "01001111",
       "01001111",
       "01001101",
       "01001011",
       "01010000",
       "01010110",
       "01010011",
       "01001100",
       "00111110",
       "00111100",
       "00110110",
       "00110000",
       "00001000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00101010",
       "00001011",
       "00111001",
       "00111001",
       "01000011",
       "01000000",
       "00111110",
       "00110110",
       "00101011",
       "00100010",
       "00001011",
       "00011010",
       "00111111",
       "01000100",
       "01001001",
       "01011011",
       "01001011",
       "01000111",
       "00101101",
       "00010010",
       "00010000",
       "00011100",
       "00010100",
       "00100110",
       "01000000",
       "01000011",
       "01000100",
       "01010010",
       "01011100",
       "01100001",
       "01011100",
       "01011011",
       "01011111",
       "01011101",
       "01011010",
       "01000110",
       "01010111",
       "01101101",
       "01011110",
       "01010001",
       "01011000",
       "01010111",
       "01010010",
       "01010010",
       "01010011",
       "01010010",
       "01010111",
       "01100000",
       "01100001",
       "01011101",
       "01011101",
       "01011010",
       "01011101",
       "01011011",
       "01010010",
       "01100010",
       "01011111",
       "01011001",
       "01000001",
       "00011101",
       "00100000",
       "00100110",
       "01010000",
       "01011000",
       "01011111",
       "01011111",
       "01100010",
       "01100100",
       "01100011",
       "01100101",
       "01101011",
       "01101111",
       "01101100",
       "01101100",
       "01101001",
       "01100111",
       "01010101",
       "01010111",
       "01010101",
       "01001111",
       "01000010",
       "01001011",
       "01011100",
       "01000101",
       "01001101",
       "01000011",
       "01001101",
       "01011100",
       "01011000",
       "01010110",
       "01011110",
       "01011001",
       "01001001",
       "01000100",
       "01000001",
       "00111111",
       "00111110",
       "00101111",
       "00001111",
       "00010000",
       "00101001",
       "01000101",
       "01000110",
       "01001110",
       "01010011",
       "01011011",
       "01011100",
       "01011101",
       "01011000",
       "01010011",
       "01010100",
       "01001001",
       "01000001",
       "00111101",
       "00110111",
       "00111010",
       "00101010",
       "00011000",
       "00000111",
       "00001011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00101111",
       "00001100",
       "00011101",
       "00100100",
       "00110011",
       "00101001",
       "00101001",
       "00100110",
       "00100100",
       "00011011",
       "00101100",
       "00100011",
       "00101111",
       "01000101",
       "01000111",
       "01011001",
       "01001101",
       "01000101",
       "00110011",
       "00010001",
       "00011010",
       "00011111",
       "00011101",
       "00110111",
       "01000110",
       "01000100",
       "01000011",
       "01001111",
       "01011101",
       "01100000",
       "01011000",
       "01011011",
       "01011110",
       "01011010",
       "01010110",
       "01011001",
       "01100000",
       "01100010",
       "01010101",
       "01001111",
       "01001111",
       "01001100",
       "01001010",
       "01001001",
       "01001001",
       "01000111",
       "01010000",
       "01100111",
       "01101100",
       "01101101",
       "01100100",
       "01010111",
       "01010110",
       "01010101",
       "01001110",
       "01011111",
       "01100010",
       "01010101",
       "01001100",
       "00100101",
       "00011110",
       "00101100",
       "01010001",
       "01010100",
       "01100001",
       "01011111",
       "01100000",
       "01011111",
       "01100000",
       "01100101",
       "01100111",
       "01100101",
       "01100110",
       "01101010",
       "01011100",
       "01010011",
       "01010000",
       "01010110",
       "01010000",
       "01010010",
       "01001101",
       "01010110",
       "01101000",
       "01100111",
       "01011101",
       "01000110",
       "01010001",
       "01011111",
       "01011101",
       "01100000",
       "01100010",
       "01011111",
       "01011010",
       "01010010",
       "01000101",
       "00111111",
       "00111110",
       "01000010",
       "00100001",
       "00001001",
       "00100101",
       "00111111",
       "01000010",
       "01001000",
       "01010010",
       "01011011",
       "01011001",
       "01010111",
       "01001100",
       "01000000",
       "00111010",
       "01000000",
       "00111110",
       "00110111",
       "00110100",
       "00101011",
       "00010110",
       "00011011",
       "00010010",
       "00011000",
       "00010001",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001111",
       "00010101",
       "00010000",
       "00011101",
       "00100000",
       "00101011",
       "00110101",
       "00111110",
       "00110110",
       "01000001",
       "00111110",
       "00111010",
       "00111011",
       "01000011",
       "01010010",
       "01011000",
       "01000010",
       "01000000",
       "00011110",
       "00101100",
       "00101000",
       "00011000",
       "01000001",
       "01000100",
       "01000011",
       "01000101",
       "01010000",
       "01011100",
       "01011100",
       "01010110",
       "01011101",
       "01100110",
       "01011001",
       "01011011",
       "01011010",
       "01010101",
       "01010011",
       "01010001",
       "01010011",
       "01001111",
       "01001011",
       "01000101",
       "01000111",
       "01000100",
       "01000000",
       "00111100",
       "01001010",
       "01011100",
       "01101111",
       "01101011",
       "01010001",
       "00111000",
       "01001110",
       "01010010",
       "01011011",
       "01011100",
       "01010010",
       "01001101",
       "00110000",
       "00011000",
       "00110111",
       "01001110",
       "01010100",
       "01100100",
       "01010101",
       "01010111",
       "01011011",
       "01100100",
       "01101010",
       "01100101",
       "01101011",
       "01101111",
       "01101110",
       "01100101",
       "01011111",
       "01010011",
       "01001110",
       "01001100",
       "01001111",
       "01010010",
       "01010101",
       "01011001",
       "01100011",
       "01100111",
       "01100110",
       "01011111",
       "01011010",
       "01011100",
       "01011011",
       "01011101",
       "01100000",
       "01011010",
       "01011010",
       "01001011",
       "01000000",
       "01000001",
       "01000010",
       "00101010",
       "00001011",
       "00010101",
       "00110100",
       "01000000",
       "01000010",
       "01010011",
       "01011001",
       "01010111",
       "01010001",
       "01000011",
       "00111110",
       "00111011",
       "00110111",
       "00110001",
       "00101101",
       "00100100",
       "00100111",
       "00101100",
       "00101110",
       "00101010",
       "00101100",
       "00011110",
       "00001011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010001",
       "00010011",
       "00010000",
       "00101011",
       "00111000",
       "00111011",
       "00111111",
       "01000101",
       "01000001",
       "00111100",
       "00111111",
       "01000110",
       "00111100",
       "01000010",
       "01010000",
       "01010111",
       "01000111",
       "01000001",
       "00110110",
       "00101100",
       "00101111",
       "00100110",
       "00110111",
       "01000010",
       "01000000",
       "01000110",
       "01010011",
       "01011101",
       "01011011",
       "01011011",
       "01011011",
       "01011111",
       "01011000",
       "01011001",
       "01001110",
       "01010000",
       "01010000",
       "01001011",
       "01001111",
       "01001010",
       "01000110",
       "01000101",
       "01001000",
       "01000101",
       "01001001",
       "01000010",
       "00101111",
       "00101010",
       "00101001",
       "00111011",
       "00101111",
       "00010111",
       "00100011",
       "00111011",
       "01010010",
       "01011001",
       "01010111",
       "01011001",
       "01001000",
       "00101001",
       "01000111",
       "01010010",
       "01010100",
       "01011001",
       "01010001",
       "01010010",
       "01011100",
       "01100011",
       "01011011",
       "01100000",
       "01110011",
       "01110101",
       "01110111",
       "01101010",
       "01000111",
       "00111010",
       "01000101",
       "01001000",
       "01000111",
       "01000111",
       "01010010",
       "01010100",
       "01010010",
       "01011010",
       "01100010",
       "01100000",
       "01011010",
       "01011110",
       "01011100",
       "01011011",
       "01100001",
       "01011011",
       "01010111",
       "01001010",
       "01000001",
       "01000000",
       "00111110",
       "00011111",
       "00010011",
       "00010011",
       "00011111",
       "01000000",
       "00111111",
       "01001000",
       "01011011",
       "01011000",
       "01001011",
       "00111100",
       "00111010",
       "00101001",
       "00011101",
       "00100010",
       "00101110",
       "00101111",
       "00111110",
       "00110000",
       "00110001",
       "00101110",
       "00110011",
       "00101000",
       "00011100",
       "00010000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010010",
       "00010001",
       "00100000",
       "01000010",
       "00111101",
       "00111111",
       "00110111",
       "00111110",
       "01000101",
       "01001001",
       "01000110",
       "01000100",
       "01000000",
       "01000001",
       "01010011",
       "01011001",
       "01010000",
       "01000010",
       "01000000",
       "00100011",
       "00011011",
       "00100000",
       "00011011",
       "01000001",
       "01000001",
       "01001000",
       "01010110",
       "01010010",
       "01010101",
       "01011100",
       "01011101",
       "01011111",
       "01011100",
       "01010010",
       "01001100",
       "01001010",
       "01001100",
       "01001011",
       "01000011",
       "01000000",
       "01000001",
       "01000110",
       "01000011",
       "01000110",
       "01000110",
       "01001010",
       "01000110",
       "00111010",
       "00011001",
       "00011000",
       "00100011",
       "00011001",
       "00011101",
       "00011110",
       "00101111",
       "01001001",
       "01010000",
       "01010110",
       "01010111",
       "01000100",
       "01011001",
       "01010111",
       "01011001",
       "01010001",
       "01010110",
       "01000111",
       "01001010",
       "01000001",
       "00110000",
       "00111101",
       "01010101",
       "01010100",
       "01010100",
       "01000010",
       "00110111",
       "01000010",
       "01000111",
       "01000110",
       "01000101",
       "01000001",
       "01001001",
       "01001011",
       "01010010",
       "01010100",
       "01010011",
       "01011111",
       "01011111",
       "01011011",
       "01011111",
       "01011100",
       "01010000",
       "01010111",
       "01011010",
       "01010011",
       "01000101",
       "00111111",
       "00110110",
       "00010100",
       "00011000",
       "00010101",
       "00010111",
       "00110010",
       "00111110",
       "01000010",
       "01011011",
       "01011100",
       "01000110",
       "00111010",
       "00101010",
       "00100011",
       "00101111",
       "00110100",
       "00111011",
       "00111010",
       "00111011",
       "00110000",
       "00111010",
       "00101010",
       "00110010",
       "00100111",
       "00101001",
       "00010101",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010110",
       "00010111",
       "00010011",
       "00110100",
       "00111101",
       "00111001",
       "01000100",
       "01000011",
       "01001100",
       "01010010",
       "01011011",
       "01010110",
       "01010110",
       "01010010",
       "01010101",
       "01011001",
       "01011110",
       "01010011",
       "01001001",
       "01000011",
       "01000000",
       "00110001",
       "00101110",
       "00110101",
       "01000100",
       "01000000",
       "01001111",
       "01010101",
       "01001111",
       "01010011",
       "01011000",
       "01100001",
       "01011010",
       "01010101",
       "01010100",
       "01001100",
       "01000100",
       "01000101",
       "01000110",
       "01000000",
       "01000011",
       "01000001",
       "01000001",
       "01000110",
       "01000011",
       "01000101",
       "01000001",
       "01000111",
       "01001010",
       "00111110",
       "00101001",
       "00100011",
       "00011100",
       "00011010",
       "00010111",
       "00011011",
       "00100110",
       "00111101",
       "00110101",
       "00100000",
       "00101000",
       "01001000",
       "01010010",
       "01010010",
       "01000000",
       "00110000",
       "00101011",
       "00101011",
       "00100011",
       "00010000",
       "00100000",
       "00100101",
       "00011111",
       "00010010",
       "00101100",
       "01001100",
       "01001110",
       "01001111",
       "01000101",
       "01000100",
       "01000000",
       "01000101",
       "01000111",
       "01001100",
       "01001110",
       "01001111",
       "01010001",
       "01010111",
       "01011010",
       "01011010",
       "01011100",
       "01010110",
       "01010110",
       "01011010",
       "01011000",
       "01001010",
       "00111101",
       "00111110",
       "00110000",
       "00100000",
       "00011100",
       "00100101",
       "00101101",
       "01000010",
       "01000110",
       "01010111",
       "01010000",
       "01000100",
       "00111000",
       "00101101",
       "00111010",
       "00111110",
       "00111000",
       "00111001",
       "00110110",
       "00111001",
       "00111101",
       "00111010",
       "00101101",
       "00101110",
       "00101001",
       "00101010",
       "00100101",
       "00010001",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010001",
       "00011010",
       "00010011",
       "00111010",
       "00111110",
       "00111100",
       "01000100",
       "01001001",
       "01001110",
       "01010100",
       "01010101",
       "01010110",
       "01011000",
       "01011011",
       "01100010",
       "01011011",
       "01011100",
       "01011010",
       "01010101",
       "01001000",
       "01000001",
       "00111111",
       "01000011",
       "01001001",
       "01000111",
       "01001101",
       "01010110",
       "01010101",
       "01010111",
       "01010100",
       "01011111",
       "01011010",
       "01010011",
       "01010001",
       "01010010",
       "01000110",
       "01001000",
       "01000100",
       "01000010",
       "01000011",
       "01000010",
       "01000000",
       "01000000",
       "01001000",
       "01000000",
       "01000011",
       "01000001",
       "01000111",
       "01000111",
       "01000101",
       "00110110",
       "00011001",
       "00011010",
       "00011001",
       "00011110",
       "00011110",
       "00011110",
       "00011111",
       "00011101",
       "00001111",
       "00010011",
       "00011010",
       "00101100",
       "00100111",
       "00011110",
       "00100100",
       "00100011",
       "00100110",
       "00011100",
       "00011000",
       "00100010",
       "00011111",
       "00011000",
       "00011101",
       "01000101",
       "01001110",
       "01001000",
       "01001110",
       "01000110",
       "01001001",
       "01001001",
       "01000101",
       "00111111",
       "01001000",
       "01000111",
       "01000111",
       "01000100",
       "01001110",
       "01010110",
       "01011000",
       "01100000",
       "01100100",
       "01011000",
       "01010111",
       "01010111",
       "01001101",
       "01000011",
       "01000011",
       "01000011",
       "00111100",
       "00110011",
       "00110011",
       "00111001",
       "01000000",
       "01000111",
       "01011101",
       "01001101",
       "01000000",
       "00110111",
       "00110111",
       "00111000",
       "00111000",
       "00111010",
       "00111101",
       "00111111",
       "01000110",
       "00111111",
       "00110010",
       "00101100",
       "00100111",
       "00101011",
       "00100111",
       "00100110",
       "00011111",
       "00100010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010001",
       "00011001",
       "00001111",
       "00101001",
       "00111101",
       "00111110",
       "00111101",
       "00111100",
       "00111110",
       "01000110",
       "00111111",
       "01000110",
       "01001011",
       "01010010",
       "01010111",
       "01011101",
       "01011010",
       "01011110",
       "01011011",
       "01010101",
       "01001001",
       "01000101",
       "01000100",
       "01001001",
       "01001111",
       "01010111",
       "01011000",
       "01011000",
       "01011011",
       "01011100",
       "01100000",
       "01010110",
       "01010011",
       "01010000",
       "01000100",
       "01000000",
       "01000010",
       "01000110",
       "01000101",
       "01000001",
       "00111110",
       "01000010",
       "00111101",
       "01000010",
       "01000111",
       "01000100",
       "01000111",
       "01001010",
       "01001010",
       "01000011",
       "00110100",
       "00011101",
       "00011101",
       "00100000",
       "00101011",
       "00110010",
       "00110111",
       "00110101",
       "00100011",
       "00011000",
       "00100001",
       "00010110",
       "00010100",
       "00010110",
       "00011000",
       "00011111",
       "00011101",
       "00101101",
       "00100110",
       "00011110",
       "00011111",
       "00011011",
       "00100001",
       "01000101",
       "01001000",
       "01000111",
       "01001001",
       "01001001",
       "01000001",
       "01000010",
       "01000111",
       "01000111",
       "01000011",
       "01000101",
       "01000100",
       "01000010",
       "01000110",
       "01010001",
       "01010110",
       "01011001",
       "01011011",
       "01011110",
       "01010111",
       "01010010",
       "01010100",
       "01010011",
       "01001101",
       "01001000",
       "00111110",
       "01000101",
       "00111110",
       "00111001",
       "00111101",
       "00111111",
       "01010001",
       "01011011",
       "01010001",
       "00111111",
       "00111001",
       "00111010",
       "00111010",
       "00111110",
       "01000100",
       "01001001",
       "01001011",
       "01001000",
       "00110100",
       "00101101",
       "00100100",
       "00100101",
       "00100111",
       "00101001",
       "00100100",
       "00101010",
       "00011110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010111",
       "00010011",
       "00010011",
       "00011011",
       "00101101",
       "00111100",
       "00111010",
       "01000001",
       "00111111",
       "00111111",
       "00111100",
       "01000010",
       "01000100",
       "01001011",
       "01010111",
       "01100000",
       "01011010",
       "01100001",
       "01100000",
       "01011101",
       "01011010",
       "01010111",
       "01010111",
       "01011100",
       "01011101",
       "01011001",
       "01011110",
       "01011011",
       "01100011",
       "01011110",
       "01011011",
       "01011101",
       "01010001",
       "01001001",
       "01000110",
       "01000001",
       "00111011",
       "01000110",
       "01001001",
       "01000000",
       "01000100",
       "01000110",
       "01000011",
       "01000011",
       "01001100",
       "01001111",
       "01001110",
       "01001011",
       "01000011",
       "00111011",
       "00100101",
       "00011101",
       "00101001",
       "00101101",
       "00110111",
       "00111001",
       "00111011",
       "00111111",
       "00111110",
       "00101011",
       "00100010",
       "00011100",
       "00100010",
       "00100000",
       "00011101",
       "00100010",
       "00011001",
       "00011101",
       "00100101",
       "00011111",
       "00011011",
       "00011001",
       "00101001",
       "01001011",
       "01000010",
       "01000111",
       "01001001",
       "01001010",
       "00111111",
       "01000010",
       "01000100",
       "01000010",
       "01000000",
       "01000101",
       "01000011",
       "01000011",
       "01000001",
       "01000010",
       "01001001",
       "01010101",
       "01010100",
       "01011110",
       "01011110",
       "01010110",
       "01010101",
       "01011000",
       "01010010",
       "01001011",
       "01001010",
       "01000101",
       "01000001",
       "00111111",
       "01000100",
       "01010011",
       "01011011",
       "01011001",
       "01010001",
       "01001011",
       "01000001",
       "01000011",
       "01000110",
       "01001001",
       "01001100",
       "01001111",
       "01001000",
       "00111011",
       "00101111",
       "00101000",
       "00100101",
       "00101100",
       "00100011",
       "00101000",
       "00100100",
       "00100111",
       "00011101",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00011010",
       "00010101",
       "00100100",
       "00101111",
       "00110110",
       "00110001",
       "00110011",
       "00110100",
       "00111000",
       "00110101",
       "00110101",
       "00111001",
       "00111010",
       "01000000",
       "00111100",
       "01001111",
       "01011110",
       "01011011",
       "01100011",
       "01011100",
       "01011111",
       "01100000",
       "01011110",
       "01100001",
       "01100100",
       "01100001",
       "01100100",
       "01100100",
       "01100001",
       "01011111",
       "01011100",
       "01011100",
       "01011000",
       "01000010",
       "00111101",
       "01000101",
       "01000000",
       "00111100",
       "01000100",
       "01001101",
       "01001000",
       "01000011",
       "01000101",
       "01000111",
       "01000110",
       "01001001",
       "01001110",
       "01010001",
       "01001101",
       "01000000",
       "00101011",
       "00100010",
       "00110110",
       "01000001",
       "00110111",
       "00111001",
       "00110000",
       "00101011",
       "00101000",
       "00111000",
       "00111010",
       "00100111",
       "00011111",
       "00011001",
       "00011101",
       "00101000",
       "00101100",
       "00100010",
       "00011111",
       "00011101",
       "00011101",
       "00010111",
       "00010100",
       "00101001",
       "01000111",
       "01000011",
       "01000110",
       "01001010",
       "01001010",
       "01000110",
       "01000101",
       "01000100",
       "00111111",
       "00111011",
       "01000101",
       "01000110",
       "01000001",
       "00111110",
       "00111001",
       "01000011",
       "01001101",
       "01010001",
       "01010111",
       "01100000",
       "01011011",
       "01011010",
       "01010101",
       "01010011",
       "01001110",
       "01010110",
       "01010010",
       "01001100",
       "01001110",
       "01010011",
       "01011110",
       "01011101",
       "01010111",
       "01010100",
       "01011010",
       "01010101",
       "01010111",
       "01011010",
       "01010110",
       "01001111",
       "01001110",
       "00111111",
       "00110011",
       "00101111",
       "00101000",
       "00101011",
       "00101011",
       "00101000",
       "00101000",
       "00100011",
       "00100101",
       "00011111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00011001",
       "00100101",
       "00111101",
       "00110110",
       "00111011",
       "00111010",
       "00111010",
       "00111000",
       "00111010",
       "00111011",
       "00110101",
       "00110011",
       "00110100",
       "00111111",
       "00111101",
       "01001100",
       "01011100",
       "01011111",
       "01011111",
       "01011111",
       "01011110",
       "01100010",
       "01011111",
       "01100011",
       "01100010",
       "01011111",
       "01100110",
       "01100100",
       "01100000",
       "01011011",
       "01011001",
       "01010000",
       "00111001",
       "00101111",
       "00110101",
       "00111011",
       "01000100",
       "01000001",
       "01000110",
       "01001001",
       "01001100",
       "01001000",
       "01001000",
       "01000111",
       "01000001",
       "00111111",
       "01001001",
       "01001001",
       "01000111",
       "01000000",
       "00110011",
       "00111100",
       "00111100",
       "00101100",
       "00101011",
       "01001000",
       "00111110",
       "00101011",
       "00101001",
       "00101111",
       "00101110",
       "00110010",
       "00100001",
       "00010100",
       "00100001",
       "00101000",
       "00011110",
       "00100000",
       "00101010",
       "00100011",
       "00011001",
       "00010111",
       "00011111",
       "00100011",
       "00111101",
       "01000110",
       "01000100",
       "01001001",
       "01001011",
       "01001010",
       "01001001",
       "01000111",
       "01000000",
       "01000001",
       "01000010",
       "01000110",
       "00111101",
       "00111100",
       "00111101",
       "01000101",
       "01000110",
       "01001001",
       "01001111",
       "01010110",
       "01010110",
       "01011011",
       "01011010",
       "01010011",
       "01010110",
       "01011011",
       "01011101",
       "01010101",
       "01011000",
       "01011001",
       "01011010",
       "01011100",
       "01011101",
       "01011010",
       "01100000",
       "01011010",
       "01010111",
       "01011001",
       "01011000",
       "01001101",
       "01001011",
       "00111010",
       "00101111",
       "00100111",
       "00101101",
       "00101010",
       "00101011",
       "00101110",
       "00101000",
       "00100011",
       "00100111",
       "00011110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001000",
       "00100010",
       "00111010",
       "00111101",
       "00111000",
       "00111100",
       "00111001",
       "00111011",
       "00111001",
       "01000001",
       "01000011",
       "01000000",
       "00111101",
       "00111101",
       "01000011",
       "01001101",
       "01011001",
       "01100011",
       "01100010",
       "01011111",
       "01100000",
       "01011100",
       "01011101",
       "01100001",
       "01100100",
       "01011111",
       "01011110",
       "01100100",
       "01100010",
       "01011101",
       "01011001",
       "01000111",
       "00101001",
       "00100011",
       "00100110",
       "00101011",
       "00111110",
       "01001100",
       "01000100",
       "01000101",
       "01000011",
       "00111101",
       "01000101",
       "01010000",
       "01001100",
       "01000001",
       "01000001",
       "01001001",
       "01000000",
       "01001001",
       "01000000",
       "00110101",
       "00110011",
       "00011110",
       "00010101",
       "00100100",
       "00111001",
       "00110101",
       "00011110",
       "00011111",
       "00100110",
       "00101100",
       "00101000",
       "00100101",
       "00101001",
       "00100011",
       "00100011",
       "00011110",
       "00010100",
       "00101101",
       "01000010",
       "00110010",
       "00011000",
       "00101000",
       "00110011",
       "00100011",
       "00111111",
       "01000101",
       "01001110",
       "01010000",
       "01001100",
       "01001001",
       "01001000",
       "01000101",
       "01000100",
       "01000101",
       "01001000",
       "01000011",
       "01000010",
       "00111111",
       "00111111",
       "01000000",
       "01000010",
       "01001000",
       "01001110",
       "01010011",
       "01010100",
       "01011010",
       "01011011",
       "01010110",
       "01011011",
       "01011101",
       "01011100",
       "01010111",
       "01011001",
       "01011100",
       "01011101",
       "01011101",
       "01011011",
       "01010111",
       "01010100",
       "01010010",
       "01010101",
       "01010110",
       "01001110",
       "01001100",
       "01000001",
       "00111001",
       "00110000",
       "00110100",
       "00110100",
       "00110111",
       "00110101",
       "00101011",
       "00100000",
       "00100010",
       "00011100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000011",
       "00010001",
       "00111000",
       "00111101",
       "00111100",
       "01000101",
       "01001000",
       "01000111",
       "01000110",
       "01001000",
       "01000101",
       "01001110",
       "01010000",
       "01010100",
       "01010011",
       "01011111",
       "01100000",
       "01011100",
       "01011111",
       "01011101",
       "01011001",
       "01011111",
       "01011011",
       "01011110",
       "01011111",
       "01011011",
       "01011101",
       "01011100",
       "01011011",
       "01011011",
       "01010110",
       "00100000",
       "00010111",
       "00100110",
       "00101001",
       "00110010",
       "01001011",
       "01001110",
       "00111101",
       "01000010",
       "00111111",
       "01000000",
       "00111100",
       "01010001",
       "01000111",
       "01000110",
       "01000101",
       "01000001",
       "01000100",
       "01000000",
       "00110000",
       "00101000",
       "00100000",
       "00010111",
       "00100010",
       "00011011",
       "00011010",
       "00100001",
       "00011010",
       "00011110",
       "00010111",
       "00100111",
       "00011001",
       "00100010",
       "00111000",
       "00110001",
       "00101011",
       "00011100",
       "00011101",
       "00100101",
       "00111000",
       "00110011",
       "00011100",
       "00010100",
       "00110101",
       "00110001",
       "00111100",
       "01000100",
       "01000110",
       "01010001",
       "01000101",
       "01000000",
       "01000100",
       "01001010",
       "01001010",
       "01000010",
       "01000111",
       "01000001",
       "01000011",
       "00111111",
       "00111100",
       "00111101",
       "01000010",
       "01000100",
       "00111111",
       "01010011",
       "01010000",
       "01010000",
       "01011100",
       "01011100",
       "01011010",
       "01010110",
       "01011101",
       "01011000",
       "01010111",
       "01011100",
       "01011110",
       "01011101",
       "01011001",
       "01010000",
       "01010010",
       "01011000",
       "01011100",
       "01011000",
       "01001110",
       "01001011",
       "01000111",
       "01000011",
       "00111101",
       "00111111",
       "00111111",
       "00111111",
       "00110011",
       "00100110",
       "00011110",
       "00100101",
       "00011010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00011101",
       "00001001",
       "00110111",
       "00111010",
       "00111110",
       "00111100",
       "01001010",
       "01001100",
       "01010011",
       "01010110",
       "01010101",
       "01011000",
       "01011011",
       "01011010",
       "01011011",
       "01010111",
       "01001101",
       "01000101",
       "01010110",
       "01011100",
       "01011100",
       "01100001",
       "01011101",
       "01011000",
       "01011100",
       "01011001",
       "01011010",
       "01011100",
       "01100000",
       "01011101",
       "01100001",
       "00100101",
       "00010100",
       "00100001",
       "00101010",
       "00110001",
       "01001111",
       "01001100",
       "01000001",
       "01000100",
       "00111111",
       "01001000",
       "00111111",
       "01001010",
       "00111111",
       "01000110",
       "00111011",
       "00111110",
       "01000001",
       "00111011",
       "00110001",
       "00101100",
       "00110001",
       "00101010",
       "00100100",
       "00011111",
       "00011111",
       "00011110",
       "00011001",
       "00100000",
       "00100110",
       "00101001",
       "00101000",
       "00100110",
       "00111110",
       "00111010",
       "00100011",
       "00011010",
       "00100001",
       "00100100",
       "00100011",
       "00011100",
       "00011010",
       "00010011",
       "00011101",
       "00110010",
       "00111101",
       "00111111",
       "00111111",
       "01000101",
       "00111101",
       "00111101",
       "00111111",
       "01001000",
       "01001000",
       "00111100",
       "01000011",
       "01000101",
       "00111100",
       "00111001",
       "00111111",
       "01000100",
       "01000111",
       "00110001",
       "00100001",
       "00110001",
       "01001000",
       "01010011",
       "01010111",
       "01011010",
       "01010101",
       "01010111",
       "01011000",
       "01011000",
       "01010111",
       "01011001",
       "01010110",
       "01010110",
       "01001011",
       "01000010",
       "01000011",
       "01000110",
       "01001011",
       "01001101",
       "01001010",
       "01001110",
       "01001000",
       "01000100",
       "01000111",
       "01000100",
       "00111011",
       "00111011",
       "00101101",
       "00101000",
       "00100000",
       "00100110",
       "00001100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000111",
       "00110000",
       "00111011",
       "00111010",
       "00110101",
       "00111110",
       "01000110",
       "01001101",
       "01000110",
       "01000101",
       "01001000",
       "01010000",
       "01010001",
       "01011000",
       "01010100",
       "01001011",
       "01001011",
       "01010111",
       "01010010",
       "01011000",
       "01011110",
       "01011100",
       "01011010",
       "01011100",
       "01011010",
       "01001110",
       "01010001",
       "01010111",
       "01011110",
       "01011111",
       "01010110",
       "00110000",
       "00100101",
       "00101101",
       "00110101",
       "01001011",
       "01000111",
       "01000000",
       "01000101",
       "01000000",
       "01000001",
       "00111110",
       "00111101",
       "00111110",
       "01000100",
       "01000010",
       "01000110",
       "01000101",
       "01001001",
       "00111100",
       "00101110",
       "00111011",
       "00101101",
       "00011011",
       "00011011",
       "00011001",
       "00011101",
       "00100001",
       "00100101",
       "00101001",
       "00101101",
       "00101111",
       "00101111",
       "00111000",
       "00110111",
       "00100000",
       "00011110",
       "00010111",
       "00100000",
       "00011001",
       "00010100",
       "00001111",
       "00010010",
       "00010010",
       "00010111",
       "00110111",
       "00111100",
       "00111100",
       "01000010",
       "01000011",
       "01001001",
       "00111100",
       "01000100",
       "01000100",
       "01000100",
       "01000011",
       "01000111",
       "01000111",
       "01000100",
       "01000111",
       "01000111",
       "01001000",
       "00101101",
       "00001101",
       "00000111",
       "00101111",
       "01010010",
       "01011001",
       "01011001",
       "01010110",
       "01010110",
       "01010010",
       "01010010",
       "01010000",
       "01010011",
       "01001110",
       "01001001",
       "00111001",
       "00111000",
       "00110000",
       "00110100",
       "00110111",
       "00111010",
       "01000001",
       "01000001",
       "00111101",
       "00111110",
       "00111011",
       "00111011",
       "00110000",
       "00110010",
       "00100100",
       "00100110",
       "00011110",
       "00101010",
       "00001000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000010",
       "00011010",
       "00111000",
       "00111000",
       "00111101",
       "00110110",
       "01000100",
       "01000000",
       "00111001",
       "00111011",
       "00111010",
       "01000011",
       "01001001",
       "01001010",
       "01010000",
       "01001011",
       "01001110",
       "01010111",
       "01001100",
       "01010110",
       "01011010",
       "01011000",
       "01010111",
       "01011000",
       "01001101",
       "00111111",
       "01000010",
       "01000011",
       "01010100",
       "01011010",
       "01011110",
       "01011011",
       "01001011",
       "01001101",
       "01010101",
       "01010110",
       "01010101",
       "01000110",
       "01000010",
       "01000100",
       "01000010",
       "01000110",
       "01000001",
       "01001000",
       "01000101",
       "01000111",
       "01000101",
       "01000100",
       "01000101",
       "00111111",
       "00110011",
       "01000010",
       "00100110",
       "00010100",
       "00011001",
       "00011101",
       "00011111",
       "00100011",
       "00100100",
       "00100111",
       "00100101",
       "00101011",
       "00101101",
       "00110100",
       "00101000",
       "00010110",
       "00100000",
       "00011101",
       "00011000",
       "00010110",
       "00010110",
       "00010011",
       "00010101",
       "00010100",
       "00011001",
       "00100101",
       "00110100",
       "00111001",
       "01000110",
       "00111000",
       "00111011",
       "00111110",
       "01000010",
       "00111111",
       "01000001",
       "00111110",
       "01000110",
       "01010101",
       "01001101",
       "01000011",
       "01000100",
       "01001000",
       "00101110",
       "00011000",
       "00011100",
       "01000010",
       "01010101",
       "01011000",
       "01011000",
       "01010101",
       "01010101",
       "01010100",
       "01001111",
       "01001100",
       "01010010",
       "01001001",
       "01000000",
       "00111011",
       "00110000",
       "00101111",
       "00110010",
       "00110010",
       "00110011",
       "00110001",
       "00110010",
       "00110011",
       "00110111",
       "00110000",
       "00101110",
       "00101010",
       "00101001",
       "00100010",
       "00100001",
       "00011110",
       "00100001",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001011",
       "00100110",
       "00110111",
       "00111011",
       "00110010",
       "00110110",
       "00110101",
       "00110101",
       "00110110",
       "00111001",
       "00111011",
       "00111110",
       "00111011",
       "00111111",
       "00111010",
       "00111100",
       "01001100",
       "01001100",
       "01010110",
       "01010100",
       "01010100",
       "01010001",
       "01010000",
       "00111100",
       "00111110",
       "00110110",
       "00111100",
       "01000110",
       "01011000",
       "01010110",
       "01010110",
       "01010110",
       "01001110",
       "01001101",
       "01001010",
       "01010101",
       "01010100",
       "01001101",
       "01000101",
       "01000000",
       "01001001",
       "01001000",
       "01001101",
       "01001011",
       "01010001",
       "01001001",
       "01000110",
       "01000101",
       "00111111",
       "00111111",
       "01000010",
       "00100100",
       "00011101",
       "00011110",
       "00100100",
       "00011111",
       "00011010",
       "00011010",
       "00100100",
       "00100110",
       "00101101",
       "00101111",
       "00111001",
       "00100011",
       "00010000",
       "00011010",
       "00011000",
       "00011011",
       "00011111",
       "00010100",
       "00010100",
       "00011011",
       "00011010",
       "00011010",
       "00010110",
       "00100010",
       "00101111",
       "00101100",
       "00100011",
       "00101111",
       "01000000",
       "01000010",
       "00111011",
       "01000001",
       "00111101",
       "01000110",
       "01001101",
       "01000100",
       "01000011",
       "01000001",
       "01001000",
       "00111101",
       "01000011",
       "01010100",
       "01011000",
       "01011001",
       "01010101",
       "01010111",
       "01010001",
       "01010010",
       "01010011",
       "01001101",
       "01001110",
       "01010110",
       "01000101",
       "00111000",
       "00111101",
       "00101000",
       "00100110",
       "00110001",
       "00101111",
       "00110011",
       "00101100",
       "00101010",
       "00110010",
       "00101111",
       "00110000",
       "00101011",
       "00100100",
       "00100110",
       "00101001",
       "00011111",
       "00100101",
       "00001100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001101",
       "00010000",
       "00101001",
       "01000000",
       "00111010",
       "00110010",
       "00111000",
       "00110111",
       "00110100",
       "00111001",
       "00110111",
       "00111011",
       "00111000",
       "00110111",
       "00111010",
       "00111100",
       "00111110",
       "00111100",
       "01010011",
       "01010100",
       "01010100",
       "01001011",
       "01000111",
       "00111011",
       "01000000",
       "00101000",
       "00110101",
       "01000000",
       "01001010",
       "01010110",
       "01010100",
       "01001001",
       "00111111",
       "00111111",
       "00111111",
       "00111111",
       "01001110",
       "01011000",
       "01001110",
       "01000111",
       "01001100",
       "01001101",
       "01010111",
       "01010001",
       "01010100",
       "01000101",
       "01000010",
       "01000001",
       "01000000",
       "01000101",
       "00101101",
       "00100100",
       "00010111",
       "00010111",
       "00100011",
       "00011101",
       "00011110",
       "00010111",
       "00011011",
       "00011111",
       "00101110",
       "00110000",
       "00111101",
       "00100110",
       "00011010",
       "00011101",
       "00011010",
       "00011111",
       "00010111",
       "00010100",
       "00010111",
       "00011010",
       "00011111",
       "00011010",
       "00011001",
       "00101010",
       "00101101",
       "00100010",
       "00101111",
       "00111110",
       "01000011",
       "01000101",
       "00111100",
       "00111010",
       "01000110",
       "01000100",
       "00111101",
       "00111011",
       "01000011",
       "01000110",
       "01010110",
       "01010110",
       "01010100",
       "01010010",
       "01010000",
       "01001111",
       "01010000",
       "01010011",
       "01010011",
       "01010100",
       "01010011",
       "01010001",
       "01010000",
       "01010100",
       "01000111",
       "00111100",
       "00111001",
       "00101101",
       "00011101",
       "00100001",
       "00101110",
       "00110100",
       "00110000",
       "00101111",
       "00110000",
       "00101101",
       "00101101",
       "00100101",
       "00100100",
       "00100001",
       "00100010",
       "00011010",
       "00100101",
       "00001010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001011",
       "00000110",
       "00101010",
       "00110101",
       "00101110",
       "00111111",
       "00101111",
       "00110101",
       "00111011",
       "00111100",
       "00111000",
       "00110001",
       "00101100",
       "00110010",
       "00111000",
       "00110101",
       "00101111",
       "01000001",
       "01010100",
       "01010101",
       "01001111",
       "01000100",
       "00111110",
       "00111110",
       "00101010",
       "00110101",
       "00111110",
       "01000100",
       "01010101",
       "01010111",
       "01000110",
       "01000000",
       "00111111",
       "00111010",
       "01000001",
       "00111101",
       "01001011",
       "01010100",
       "01011011",
       "01011010",
       "01010110",
       "01011010",
       "01001010",
       "01000001",
       "00111111",
       "00111100",
       "00111010",
       "01000110",
       "00110111",
       "00100101",
       "00100100",
       "00011011",
       "00011110",
       "00011110",
       "00011000",
       "00011010",
       "00011000",
       "00011000",
       "00011000",
       "00100110",
       "00101010",
       "00110011",
       "00100000",
       "00010010",
       "00100001",
       "00100011",
       "00100101",
       "00011100",
       "00100000",
       "00011011",
       "00011010",
       "00011111",
       "00011101",
       "00100110",
       "00110001",
       "00110110",
       "00101101",
       "00111110",
       "01000000",
       "00111111",
       "01000100",
       "01000010",
       "00111111",
       "01000110",
       "01000101",
       "00111110",
       "00111111",
       "01000101",
       "01001101",
       "01010011",
       "01001010",
       "01000010",
       "01000100",
       "01001001",
       "01010000",
       "01010010",
       "01010101",
       "01010000",
       "01001011",
       "01001110",
       "01010010",
       "01010001",
       "01010110",
       "01001001",
       "00111101",
       "00110110",
       "00101101",
       "00011111",
       "00010110",
       "00100000",
       "00110010",
       "00110000",
       "00110100",
       "00101100",
       "00101011",
       "00101010",
       "00100100",
       "00100110",
       "00100101",
       "00011011",
       "00100001",
       "00011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000100",
       "00011001",
       "00101000",
       "00011011",
       "00100101",
       "00110010",
       "00111011",
       "00111001",
       "00110001",
       "00101100",
       "00100110",
       "00100101",
       "00101101",
       "00110011",
       "00110010",
       "00111100",
       "01001011",
       "01001101",
       "01001100",
       "01000100",
       "00111110",
       "00111111",
       "00101110",
       "00111010",
       "00111101",
       "01000011",
       "01010010",
       "01010110",
       "01001001",
       "01000001",
       "01000010",
       "00101101",
       "00111100",
       "00111010",
       "01000010",
       "01001011",
       "01010110",
       "01011000",
       "01010100",
       "01001011",
       "00111110",
       "01000011",
       "00111100",
       "00111001",
       "00111110",
       "00110101",
       "00011100",
       "00011111",
       "00100000",
       "00100011",
       "00100100",
       "00011100",
       "00011100",
       "00011000",
       "00011010",
       "00010111",
       "00011100",
       "00100101",
       "00101000",
       "00110000",
       "00011001",
       "00001111",
       "00011001",
       "00011001",
       "00011110",
       "00011010",
       "00011001",
       "00010100",
       "00010111",
       "00010111",
       "00100001",
       "00101011",
       "00101110",
       "00111010",
       "00101111",
       "00111010",
       "01000000",
       "01000010",
       "01000101",
       "01000111",
       "01001011",
       "01000101",
       "01001001",
       "01000101",
       "01000100",
       "01001100",
       "01001110",
       "01000010",
       "01000000",
       "00111010",
       "00111100",
       "00111011",
       "01001011",
       "01010100",
       "01010110",
       "01001011",
       "00111001",
       "00111100",
       "01001101",
       "01010000",
       "01010100",
       "01001101",
       "01000001",
       "00111001",
       "00110001",
       "00100011",
       "00100001",
       "00010000",
       "00100000",
       "00101111",
       "00110110",
       "00110001",
       "00101001",
       "00100100",
       "00101010",
       "00101010",
       "00100100",
       "00010110",
       "00100011",
       "00001011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000010",
       "00001011",
       "00001101",
       "00100011",
       "00101001",
       "00101111",
       "00101010",
       "00101010",
       "00101100",
       "00110011",
       "00101000",
       "00101110",
       "00110101",
       "00110011",
       "00111100",
       "01000001",
       "01001011",
       "01001001",
       "00111101",
       "00111001",
       "00111101",
       "00101110",
       "00110010",
       "01000001",
       "00111111",
       "01001110",
       "01010101",
       "01001100",
       "01000000",
       "01000010",
       "00110110",
       "00110000",
       "00111010",
       "00111101",
       "01000001",
       "01000100",
       "01000101",
       "01000011",
       "00111100",
       "01000000",
       "00111001",
       "00110011",
       "00111000",
       "00111010",
       "00100001",
       "00010110",
       "00011010",
       "00100000",
       "00011110",
       "00100010",
       "00100100",
       "00011100",
       "00010111",
       "00011001",
       "00011010",
       "00011001",
       "00100011",
       "00101010",
       "00110000",
       "00011000",
       "00001111",
       "00010011",
       "00011001",
       "00011010",
       "00010101",
       "00010001",
       "00010101",
       "00011000",
       "00001111",
       "00011001",
       "00011010",
       "00010010",
       "00110111",
       "00110001",
       "00110111",
       "01000001",
       "00111110",
       "01001011",
       "01001010",
       "01001001",
       "01000000",
       "01001000",
       "01000101",
       "01001011",
       "01001111",
       "01001000",
       "00111010",
       "00111010",
       "00110111",
       "00110111",
       "00111000",
       "01001001",
       "01001111",
       "01010000",
       "01000011",
       "00110111",
       "00110101",
       "01000101",
       "01010101",
       "01010010",
       "01001111",
       "01001001",
       "00111000",
       "00111000",
       "00110000",
       "00110010",
       "00100000",
       "00010110",
       "00011111",
       "00101111",
       "00110010",
       "00101111",
       "00100111",
       "00100111",
       "00011111",
       "00011000",
       "00011000",
       "00001110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010010",
       "00000101",
       "00010010",
       "00011010",
       "00011010",
       "00100100",
       "00101101",
       "00101111",
       "00110110",
       "00110010",
       "00110100",
       "00110011",
       "00110000",
       "00111001",
       "00110111",
       "01000001",
       "01001000",
       "00111100",
       "00111001",
       "00111100",
       "00110011",
       "00101100",
       "00111100",
       "00111100",
       "01001001",
       "01010011",
       "01001010",
       "01000100",
       "00111111",
       "00111101",
       "00101110",
       "00110001",
       "01000001",
       "00111110",
       "00111111",
       "00111111",
       "01000000",
       "01000010",
       "01000010",
       "00110111",
       "01000101",
       "01000011",
       "01000110",
       "00111000",
       "00100001",
       "00011101",
       "00011001",
       "00011010",
       "00100010",
       "00011011",
       "00011111",
       "00011000",
       "00011001",
       "00010100",
       "00010111",
       "00101000",
       "00100110",
       "00110000",
       "00100011",
       "00010011",
       "00010001",
       "00010101",
       "00010011",
       "00010100",
       "00010110",
       "00010110",
       "00010110",
       "00001100",
       "00010011",
       "00010111",
       "00010000",
       "00101001",
       "00111000",
       "00101111",
       "00111101",
       "00111100",
       "01000101",
       "01010001",
       "01010101",
       "01001011",
       "01001100",
       "01010000",
       "01010011",
       "01000100",
       "00111100",
       "00111100",
       "00110110",
       "00110101",
       "00111111",
       "00111100",
       "01001101",
       "01010011",
       "01001010",
       "00110101",
       "00110001",
       "00110001",
       "00111000",
       "01010000",
       "01010011",
       "01010010",
       "01010001",
       "00111110",
       "00110111",
       "00110001",
       "00111000",
       "00110100",
       "00101010",
       "00011100",
       "00011100",
       "00011011",
       "00011111",
       "00011101",
       "00010100",
       "00010100",
       "00010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001101",
       "00001101",
       "00011011",
       "00011001",
       "00101011",
       "00101111",
       "00110001",
       "00101011",
       "00110110",
       "00110010",
       "00110110",
       "00110001",
       "00110011",
       "00110010",
       "00110101",
       "01001101",
       "01000001",
       "00110100",
       "00111000",
       "00111101",
       "00110101",
       "00110101",
       "01000010",
       "00111110",
       "01001011",
       "01001101",
       "01001100",
       "00111110",
       "00111100",
       "00110111",
       "00101101",
       "00110101",
       "00111010",
       "00111011",
       "01000001",
       "00111001",
       "00110010",
       "00100100",
       "00111001",
       "01001101",
       "01001011",
       "01001101",
       "01000101",
       "00101001",
       "00011001",
       "00010011",
       "00011000",
       "00011101",
       "00011011",
       "00011010",
       "00011100",
       "00010111",
       "00010101",
       "00011001",
       "00100100",
       "00100011",
       "00100111",
       "00100100",
       "00010110",
       "00010000",
       "00001010",
       "00010010",
       "00011010",
       "00010111",
       "00010000",
       "00010001",
       "00001110",
       "00001110",
       "00010010",
       "00010011",
       "00011111",
       "00111010",
       "00110110",
       "00110101",
       "01000010",
       "01000000",
       "01001011",
       "01010100",
       "01011001",
       "01010010",
       "01001111",
       "01000101",
       "01000001",
       "00111111",
       "00110011",
       "00101110",
       "01000000",
       "00111111",
       "00111111",
       "01001000",
       "01010010",
       "01000000",
       "00110010",
       "00101010",
       "00101111",
       "00110011",
       "01000110",
       "01010010",
       "01010010",
       "01010100",
       "01000111",
       "00111110",
       "00110110",
       "00110001",
       "00110011",
       "00110011",
       "00110001",
       "00100110",
       "00011010",
       "00001101",
       "00010001",
       "00001000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001001",
       "00000100",
       "00100001",
       "00011101",
       "00101111",
       "00110001",
       "00110101",
       "00110010",
       "00111000",
       "00110010",
       "00110100",
       "00110011",
       "00110001",
       "00110110",
       "00110101",
       "01001010",
       "01000110",
       "00111110",
       "00110101",
       "00110101",
       "00111010",
       "00111011",
       "01000000",
       "00111010",
       "01000000",
       "01001001",
       "01001010",
       "01000000",
       "00111010",
       "00111111",
       "00101101",
       "00100011",
       "00101110",
       "00101100",
       "00100100",
       "00011111",
       "00010100",
       "00001111",
       "00001010",
       "00101000",
       "00101111",
       "00110011",
       "00111000",
       "00101111",
       "00100101",
       "00011101",
       "00011001",
       "00010011",
       "00011000",
       "00010111",
       "00011010",
       "00011001",
       "00100010",
       "00011001",
       "00100011",
       "00011011",
       "00011110",
       "00100101",
       "00011001",
       "00010011",
       "00001101",
       "00010100",
       "00100000",
       "00010111",
       "00010010",
       "00001101",
       "00010011",
       "00001100",
       "00001110",
       "00010000",
       "00010001",
       "00011001",
       "00101010",
       "00110010",
       "00111101",
       "00111110",
       "00111101",
       "01000101",
       "01001110",
       "01001101",
       "01001000",
       "00111000",
       "00111110",
       "00110110",
       "00101000",
       "00110011",
       "00111111",
       "00111001",
       "01000001",
       "01001110",
       "01001011",
       "00111011",
       "00110101",
       "00101111",
       "00110000",
       "00111000",
       "01000001",
       "01010001",
       "01010000",
       "01010100",
       "01010000",
       "01001010",
       "01000010",
       "00111010",
       "00110100",
       "00110010",
       "00110001",
       "00110001",
       "00101001",
       "00011110",
       "00001000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010100",
       "00000100",
       "00010101",
       "00011011",
       "00100011",
       "00101010",
       "00110011",
       "00110011",
       "00100101",
       "00011111",
       "00100110",
       "00101110",
       "00101101",
       "00101100",
       "00101010",
       "00110111",
       "01000101",
       "01010110",
       "01001011",
       "00110101",
       "00111010",
       "00111110",
       "00111100",
       "01000000",
       "01000010",
       "01000010",
       "00111111",
       "00111111",
       "00111001",
       "00110111",
       "00111100",
       "00100100",
       "00011100",
       "00001110",
       "00010100",
       "00011011",
       "00011101",
       "00100001",
       "00011100",
       "00001010",
       "00010000",
       "00010111",
       "00110000",
       "00111100",
       "00110010",
       "00101000",
       "00011100",
       "00010111",
       "00010101",
       "00011100",
       "00011100",
       "00011111",
       "00011111",
       "00011001",
       "00101000",
       "00011110",
       "00100010",
       "00100100",
       "00100101",
       "00010110",
       "00011001",
       "00010110",
       "00011101",
       "00011001",
       "00010000",
       "00001011",
       "00010011",
       "00010100",
       "00011111",
       "00010101",
       "00010110",
       "00100100",
       "00100110",
       "00101111",
       "00101101",
       "00110101",
       "00110111",
       "00111011",
       "01000001",
       "01000110",
       "01000011",
       "00111011",
       "00111000",
       "00011111",
       "00101101",
       "00111010",
       "00110101",
       "00111100",
       "01000011",
       "01001101",
       "01000001",
       "00111101",
       "00110110",
       "00101110",
       "00101101",
       "00111001",
       "00111011",
       "01001110",
       "01001011",
       "01010001",
       "01001111",
       "01001000",
       "01001010",
       "01001110",
       "00111110",
       "00111010",
       "00101110",
       "00110010",
       "00101001",
       "00101100",
       "00010000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001100",
       "00000011",
       "00001110",
       "00010001",
       "00011110",
       "00100110",
       "00110001",
       "00010010",
       "00100101",
       "00100101",
       "00110111",
       "00110000",
       "00101010",
       "00101110",
       "00110001",
       "00111000",
       "01000101",
       "01001101",
       "01000101",
       "00111100",
       "01000000",
       "00111110",
       "00111100",
       "01000011",
       "01000001",
       "00111100",
       "00111010",
       "00111001",
       "00111101",
       "00110011",
       "00010001",
       "00000111",
       "00001010",
       "00010110",
       "00011110",
       "00011111",
       "00011101",
       "00100100",
       "00011110",
       "00001011",
       "00001110",
       "00000000",
       "00111101",
       "00111001",
       "00101111",
       "00100010",
       "00011110",
       "00010111",
       "00100000",
       "00100010",
       "00100001",
       "00011100",
       "00011101",
       "00011110",
       "00011011",
       "00100101",
       "00011110",
       "00100100",
       "00010101",
       "00011000",
       "00010110",
       "00011000",
       "00010110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00110000",
       "00100110",
       "00111010",
       "00111101",
       "00110110",
       "00101100",
       "00101110",
       "00110101",
       "00111011",
       "00110111",
       "00111100",
       "00110111",
       "00111100",
       "00101111",
       "00100101",
       "00111010",
       "00110111",
       "00110110",
       "00111111",
       "01000111",
       "00111111",
       "00111001",
       "00111001",
       "00110100",
       "00100000",
       "00110000",
       "00110110",
       "00111010",
       "01001001",
       "01000010",
       "01001011",
       "01000011",
       "01000101",
       "01000101",
       "01001111",
       "01000111",
       "01000100",
       "00110000",
       "00101101",
       "00100100",
       "00101110",
       "00011010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001001",
       "00000101",
       "00001010",
       "00010010",
       "00100101",
       "00001100",
       "00010001",
       "00001110",
       "00011010",
       "00101010",
       "00110000",
       "00101111",
       "00110010",
       "00101100",
       "00110011",
       "00110100",
       "00111101",
       "01000100",
       "01000010",
       "01000100",
       "00111010",
       "00111000",
       "01000011",
       "00111110",
       "01000010",
       "00111100",
       "00110101",
       "00011111",
       "00001110",
       "00001101",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00111010",
       "00110011",
       "00100001",
       "00011011",
       "00011000",
       "00011010",
       "00011110",
       "00011010",
       "00011011",
       "00100010",
       "00100100",
       "00011010",
       "00101100",
       "00100010",
       "00100011",
       "00010001",
       "00011101",
       "00010011",
       "00001111",
       "00001110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00111000",
       "00110001",
       "00110100",
       "00111001",
       "00111111",
       "01001001",
       "00111100",
       "00110001",
       "00111111",
       "00111100",
       "00111001",
       "00111000",
       "00110101",
       "00100001",
       "00110011",
       "00110101",
       "00111010",
       "01000010",
       "01000101",
       "00111101",
       "00111000",
       "00110011",
       "00110011",
       "00101010",
       "00100111",
       "00110101",
       "00111000",
       "01000000",
       "00111111",
       "00111110",
       "00111010",
       "00110101",
       "00111001",
       "00110110",
       "00111111",
       "01000010",
       "01000010",
       "00110001",
       "00101100",
       "00100100",
       "00101101",
       "00011100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000111",
       "00001000",
       "00000101",
       "00001000",
       "00000110",
       "00001100",
       "00001100",
       "00000111",
       "00011010",
       "00100100",
       "00110010",
       "00110001",
       "00110010",
       "00110000",
       "00110000",
       "00111010",
       "00111110",
       "00111100",
       "00110000",
       "00100101",
       "00111100",
       "00110100",
       "00101000",
       "00011110",
       "00010010",
       "00001010",
       "00000111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00110111",
       "00101010",
       "00011101",
       "00010011",
       "00010110",
       "00001110",
       "00010110",
       "00010111",
       "00011010",
       "00011100",
       "00100010",
       "00011110",
       "00101100",
       "00101101",
       "00100101",
       "00011100",
       "00011101",
       "00010111",
       "00001110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00100001",
       "00101001",
       "00110000",
       "00011111",
       "00110000",
       "00111011",
       "00111010",
       "00101100",
       "00110000",
       "00110001",
       "00110100",
       "00101001",
       "00011101",
       "00101111",
       "00111100",
       "00110101",
       "00111001",
       "00111110",
       "00111111",
       "00110111",
       "00110111",
       "00110011",
       "00110010",
       "00101010",
       "00111000",
       "00110010",
       "00111000",
       "00111100",
       "00111110",
       "00110111",
       "00101101",
       "00101110",
       "00101011",
       "00101010",
       "00111000",
       "00110111",
       "00110100",
       "00110001",
       "00101001",
       "00100011",
       "00101010",
       "00011100",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000111",
       "00001000",
       "00001110",
       "00100011",
       "00110010",
       "00101000",
       "00100110",
       "00100100",
       "00101010",
       "00100100",
       "00011001",
       "00011001",
       "00010111",
       "00011101",
       "00001111",
       "00001101",
       "00001001",
       "00001101",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00100110",
       "00100000",
       "00011100",
       "00010101",
       "00000000",
       "00011001",
       "00011010",
       "00011011",
       "00010110",
       "00011001",
       "00011111",
       "00100100",
       "00101001",
       "00011111",
       "00011111",
       "00010110",
       "00010110",
       "00010000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010011",
       "00010101",
       "00001111",
       "00010011",
       "00001010",
       "00001101",
       "00001101",
       "00010110",
       "00101000",
       "00100111",
       "00100110",
       "00011010",
       "00101101",
       "00110111",
       "00110110",
       "00110110",
       "00110100",
       "00110111",
       "00110111",
       "00110101",
       "00110000",
       "00101110",
       "00110011",
       "00110011",
       "00101101",
       "00111010",
       "00111001",
       "00111011",
       "00110011",
       "00101011",
       "00101100",
       "00101010",
       "00101001",
       "00101101",
       "00110001",
       "00101011",
       "00101100",
       "00100001",
       "00101011",
       "00100101",
       "00011010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001100",
       "00001101",
       "00010100",
       "00011110",
       "00010101",
       "00010110",
       "00010001",
       "00011001",
       "00100000",
       "00010111",
       "00000111",
       "00001111",
       "00001010",
       "00001101",
       "00010011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010001",
       "00001110",
       "00010011",
       "00010111",
       "00011110",
       "00010101",
       "00100011",
       "00100100",
       "00011001",
       "00010111",
       "00010101",
       "00010011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001111",
       "00010110",
       "00010111",
       "00010110",
       "00001101",
       "00001111",
       "00001001",
       "00001010",
       "00011011",
       "00011000",
       "00011100",
       "00100010",
       "00101001",
       "00110101",
       "00110000",
       "00110100",
       "00101110",
       "00110000",
       "00101111",
       "00101111",
       "00101011",
       "00110110",
       "00110100",
       "00110000",
       "00110011",
       "00111011",
       "00110011",
       "00110000",
       "00101010",
       "00101010",
       "00101100",
       "00101000",
       "00101000",
       "00100111",
       "00101010",
       "00100111",
       "00101101",
       "00100111",
       "00100011",
       "00100010",
       "00001111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001010",
       "00010001",
       "00001011",
       "00010010",
       "00001100",
       "00001010",
       "00001010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010100",
       "00010110",
       "00100001",
       "00011111",
       "00100110",
       "00101010",
       "00011100",
       "00010110",
       "00010010",
       "00010101",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00011001",
       "00000000",
       "00000000",
       "00010011",
       "00011101",
       "00001110",
       "00010011",
       "00010101",
       "00011101",
       "00101110",
       "00110111",
       "00110100",
       "00101110",
       "00100111",
       "00100111",
       "00101000",
       "00110001",
       "00110101",
       "00110011",
       "00110101",
       "00110110",
       "00110000",
       "00101001",
       "00101110",
       "00101011",
       "00101000",
       "00101001",
       "00100101",
       "00100110",
       "00100111",
       "00101001",
       "00101110",
       "00100111",
       "00100100",
       "00010111",
       "00100000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010010",
       "00010010",
       "00010100",
       "00011011",
       "00100001",
       "00011111",
       "00010100",
       "00001010",
       "00001101",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000101",
       "00001010",
       "00000111",
       "00001001",
       "00010011",
       "00011111",
       "00011111",
       "00011010",
       "00101001",
       "00110111",
       "00111001",
       "00110000",
       "00110011",
       "00101111",
       "00101101",
       "00101010",
       "00101111",
       "00101011",
       "00101110",
       "00100111",
       "00011111",
       "00011100",
       "00100001",
       "00011111",
       "00011110",
       "00011110",
       "00010110",
       "00001111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010000",
       "00010010",
       "00011000",
       "00011111",
       "00011100",
       "00010000",
       "00001001",
       "00010101",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001101",
       "00001011",
       "00001110",
       "00010011",
       "00011100",
       "00011011",
       "00110010",
       "00111101",
       "00110010",
       "00110000",
       "00101000",
       "00101000",
       "00101001",
       "00101011",
       "00100111",
       "00100101",
       "00011101",
       "00010010",
       "00000111",
       "00010011",
       "00001101",
       "00001110",
       "00001010",
       "00000110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00011000",
       "00010101",
       "00010111",
       "00011000",
       "00011010",
       "00001111",
       "00010000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00011000",
       "00011111",
       "00101110",
       "00111100",
       "00101101",
       "00101010",
       "00101010",
       "00101000",
       "00100101",
       "00011011",
       "00010101",
       "00001100",
       "00001111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00010011",
       "00010010",
       "00010111",
       "00011000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00100100",
       "00100010",
       "00011100",
       "00011101",
       "00100000",
       "00010101",
       "00001000",
       "00010000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00001011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000"
        );

begin

  addr1_int <= TO_INTEGER(unsigned(addr1));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout1 <= filaimg(addr1_int);
    end if;
  end process;

end BEHAVIORAL;
